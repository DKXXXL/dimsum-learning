From dimsum.core Require Export module trefines.
From dimsum.core.iris Require Export sat sim expr combinators.

(** This file reexports all relevant modules and should be imported by clients. *)
