Require Import refframe.base.
Require Import stdpp.namespaces.
Require Import stdpp.strings.
Require Import stdpp.gmap.
Require Import stdpp.binders.
Require Import stdpp.propset.

Inductive event (EV : Type) : Type :=
| Ub | Vis (e : EV).
Arguments Ub {_}.
Arguments Vis {_}.

(*** angelic module *)
Record module (EV : Type) : Type := {
  m_state : Type;
  m_step : m_state → option EV → (m_state → Prop) → Prop;
  (* TODO: we probably want to add the following:
-  m_step_proper σ κ : Proper ((pointwise_relation m_state impl) ==> impl) (m_step σ κ);
*)
}.

Arguments m_state {_}.
Arguments m_step {_}.

Inductive has_trace {EV} (m : module EV) : m.(m_state) → list (event EV) → (m.(m_state) → Prop) → Prop :=
| TraceEnd σ (Pσ : _ → Prop):
    Pσ σ →
    has_trace m σ [] Pσ
| TraceStep σ1 Pσ2 Pσ3 κ κs:
    m.(m_step) σ1 κ Pσ2 →
    (∀ σ2, Pσ2 σ2 → has_trace m σ2 κs Pσ3) →
    has_trace m σ1 (option_list (Vis <$> κ) ++ κs) Pσ3
.
Notation " σ '~{' m , κ '}~>' σ' " := (has_trace m σ κ σ') (at level 40).

Global Instance has_trace_proper {EV} (m : module EV) :
  Proper ((=) ==> (=) ==> (pointwise_relation m.(m_state) impl) ==> impl) (has_trace m).
Proof.
  move => ?? -> ?? -> Pσ1 Pσ2 HP Ht.
  elim: Ht Pσ2 HP.
  - move => ???? HP. apply: TraceEnd. by apply: HP.
  - move => ??????????. apply: TraceStep; naive_solver.
Qed.

(* This should capture that the events on the trace don't depend on
angelic choices. This is currently a precondition for horizontal
compositionality. TODO: Is this really necessary? *)
Definition angelic_trace_det {EV} (m : module EV) : Prop :=
  (∀ σ1 e Pσ1, m_step m σ1 e Pσ1 → (¬ ∃ σ, Pσ1 σ) ∨ ∃ σ, Pσ1 σ ∧ (∀ κs σ3, Pσ1 σ3 → σ ~{ m, κs }~> (λ _, True) → σ3 ~{ m, κs }~> (λ _, True))).

Lemma TraceStep' {EV} κs κs' (m : module EV) Pσ2 σ1 Pσ3 κ :
  m.(m_step) σ1 κ Pσ2 →
  κs = option_list (Vis <$> κ) ++ κs' →
  (∀ σ2, Pσ2 σ2 → σ2 ~{ m, κs' }~> Pσ3) →
  σ1 ~{ m, κs }~> Pσ3.
Proof. move => ? -> ?. by apply: TraceStep. Qed.

Lemma has_trace_trans {EV} κs1 κs2 (m : module EV) σ1 Pσ2 σ3 :
  σ1 ~{ m, κs1 }~> Pσ2 →
  (∀ σ2, Pσ2 σ2 → σ2 ~{ m, κs2 }~> σ3) →
  σ1 ~{ m, κs1 ++ κs2 }~> σ3.
Proof.
  elim; eauto.
  move => ?????????. rewrite -app_assoc. econstructor; eauto.
Qed.

Lemma has_trace_add_empty {EV} κs1 (m : module EV) σ1 Pσ2:
  σ1 ~{ m, κs1 ++ [] }~> Pσ2 →
  σ1 ~{ m, κs1 }~> Pσ2.
Proof. by rewrite -{2}[κs1](right_id_L [] (++)). Qed.

Lemma has_trace_ub_inv {EV} κs (m : module EV) σ1 Pσ1':
  σ1 ~{m, Ub :: κs }~> Pσ1' →
  σ1 ~{ m, [] }~> (λ σ3, False).
Proof.
  move Hκ: (Ub :: κs) => κ Hκs.
  elim: Hκs Hκ => //.
  move => ??? [] //= ??? IH ?.
  apply: TraceStep' => //. naive_solver.
Qed.

Lemma has_trace_cons_inv {EV} κs κ (m : module EV) σ1 Pσ3:
  σ1 ~{ m, Vis κ :: κs }~> Pσ3 →
  σ1 ~{ m, [] }~> (λ σ2, ∃ Pσ, m.(m_step) σ2 (Some κ) Pσ ∧ (∀ σ2', Pσ σ2' → σ2' ~{ m, κs }~> Pσ3)).
Proof.
  move Hs: (Vis κ :: κs) => s Hκs.
  elim: Hκs Hs => //.
  move => ??? [] //=.
  + move => ???? IH [] ??. subst. apply: TraceEnd. eexists _. by split.
  + move => ??? IH ?. apply: TraceStep' => //. naive_solver.
Qed.

Lemma has_trace_app_inv {EV} κs1 κs2 (m : module EV) σ1 σ3:
  σ1 ~{ m, κs1 ++ κs2 }~> σ3 →
  σ1 ~{ m, κs1 }~> (λ σ2, σ2 ~{ m, κs2 }~> σ3).
Proof.
  elim: κs1 σ1 => /=. { move => ??. by apply: TraceEnd. }
  move => [|?] ? IH ?.
  - move => /has_trace_ub_inv ?. by apply: (has_trace_trans []).
  - move => /(has_trace_cons_inv _ _)?.
    apply: (has_trace_trans []) => //= ?[?[??]].
    apply: TraceStep'; [done..|]. naive_solver.
Qed.

Lemma has_trace_ub_app_inv {EV} κs (m : module EV) σ1 σ2:
  σ1 ~{ m, κs ++ [Ub] }~> σ2 → σ1 ~{ m, κs }~> (λ _, False).
Proof.
  move => /has_trace_app_inv?.
  apply: has_trace_add_empty.
  apply: has_trace_trans; [done|] => /= ??.
  by apply: has_trace_ub_inv.
Qed.

Record mod_state EV := MS {
  ms_module : module EV;
  ms_state : ms_module.(m_state);
}.
Arguments MS {_}.
Arguments ms_module {_}.
Arguments ms_state {_}.
Coercion ms_module : mod_state >-> module.

Record refines {EV} (mimpl mspec : mod_state EV) : Prop := {
  ref_subset:
    ∀ κs, mimpl.(ms_state) ~{ mimpl, κs }~> (λ _, True) → mspec.(ms_state) ~{ mspec, κs }~> (λ _, True)
}.

Global Instance sqsubseteq_refines EV : SqSubsetEq (mod_state EV) := refines.

Definition refines_equiv {EV} (m1 m2 : mod_state EV) : Prop := m1 ⊑ m2 ∧ m2 ⊑ m1.

Global Instance equiv_refines EV : Equiv (mod_state EV) := refines_equiv.


(*** demonic module with only degenerate angelic non-determinism *)

Record dem_module (EV : Type) : Type := {
  dm_state : Type;
  dm_step : dm_state → option EV → dm_state → Prop;
  dm_is_ub : dm_state → Prop;
}.
Arguments dm_state {_}.
Arguments dm_step {_}.
Arguments dm_is_ub {_}.

Inductive dem_has_trace {EV} (m : dem_module EV) : m.(dm_state) → list (event EV) → m.(dm_state) → Prop :=
| DemTraceEnd σ:
    dem_has_trace m σ [] σ
| DemTraceStep σ1 σ2 σ3 κ κs:
    m.(dm_step) σ1 κ σ2 →
    dem_has_trace m σ2 κs σ3 →
    dem_has_trace m σ1 (option_list (Vis <$> κ) ++ κs) σ3
| DemTraceUb σ1 κs σ2:
    m.(dm_is_ub) σ1 →
    dem_has_trace m σ1 κs σ2
.
Notation " σ '~{' m , κ '}~>ₘ' σ' " := (dem_has_trace m σ κ σ') (at level 40).
Notation " σ '~{' m , κ '}~>ₘ' - " := (∃ σ', dem_has_trace m σ κ σ') (at level 40).

Lemma DemTraceStep' {EV} κs κs' (m : dem_module EV) σ2 σ1 σ3 κ :
  m.(dm_step) σ1 κ σ2 →
  κs = option_list (Vis <$> κ) ++ κs' →
  σ2 ~{ m, κs' }~>ₘ σ3 →
  σ1 ~{ m, κs }~>ₘ σ3.
Proof. move => ? -> ?. by apply: DemTraceStep. Qed.

Lemma DemTraceUbRefl {EV} (m : dem_module EV) σ κs :
  m.(dm_is_ub) σ →
  σ ~{ m, κs }~>ₘ σ.
Proof. move => ?. by apply: DemTraceUb. Qed.

Lemma dem_has_trace_trans {EV} κs1 κs2 (m : dem_module EV) σ1 σ2 σ3 :
  σ1 ~{ m, κs1 }~>ₘ σ2 →
  σ2 ~{ m, κs2 }~>ₘ σ3 →
  σ1 ~{ m, κs1 ++ κs2 }~>ₘ σ3.
Proof.
  elim => //.
  - move => ?????????. rewrite -app_assoc. econstructor; eauto.
  - move => ?????. by apply: DemTraceUb.
Qed.

Lemma dem_has_trace_add_empty {EV} κs1 (m : dem_module EV) σ1 σ2 :
  σ1 ~{ m, κs1 ++ [] }~>ₘ σ2 →
  σ1 ~{ m, κs1 }~>ₘ σ2.
Proof. by rewrite -{2}[κs1](right_id_L [] (++)). Qed.

Lemma dem_has_trace_ub_inv {EV} κs (m : dem_module EV) σ1 σ2:
  σ1 ~{m, Ub :: κs }~>ₘ σ2 →
  ∃ σ3, σ1 ~{ m, [] }~>ₘ σ3 ∧ m.(dm_is_ub) σ3.
Proof.
  move Hκ: (Ub :: κs) => κ Hκs.
  elim: Hκs Hκ => //.
  - move => ??? [] //= ??? IH ?. have [//|?[??]]:= IH.
    eexists _. split => //. by apply: DemTraceStep'.
  - move => ?????. eexists. split => //. by apply: DemTraceUb.
Qed.

Lemma dem_has_trace_cons_inv {EV} κs κ (m : dem_module EV) σ1 σ3:
  σ1 ~{ m, Vis κ :: κs }~>ₘ σ3 →
  ∃ σ2 σ2', σ1 ~{ m, [] }~>ₘ σ2 ∧ (m.(dm_is_ub) σ2 ∨ m.(dm_step) σ2 (Some κ) σ2' ∧ σ2' ~{ m, κs }~>ₘ σ3).
Proof.
  move Hs: (Vis κ :: κs) => s Hκs.
  elim: Hκs Hs => //.
  - move => ??? [] //=.
    + move => ???? IH [] ??. subst. eexists _, _. split. by apply DemTraceEnd. right. naive_solver.
    + move => ??? IH ?. have [//|?[?[??]]]:= IH. eexists _, _. split; [ | done]. by apply: DemTraceStep'.
  - move => ?????. eexists _, σ1. split; [ | by left]. by apply: DemTraceEnd.
Qed.

Lemma dem_has_trace_app_inv {EV} κs1 κs2 (m : dem_module EV) σ1 σ3:
  σ1 ~{ m, κs1 ++ κs2 }~>ₘ σ3 →
  ∃ σ2, σ1 ~{ m, κs1 }~>ₘ σ2 ∧ σ2 ~{ m, κs2 }~>ₘ σ3.
Proof.
  elim: κs1 σ1 => /=. { move => ?. eexists. split => //. apply: DemTraceEnd. }
  move => [|?] ? IH ?.
  - move => /dem_has_trace_ub_inv[σ' [??]]. eexists σ'. split; [| by apply DemTraceUb].
    apply: (dem_has_trace_trans []) => //. by apply DemTraceUb.
  - move => /(dem_has_trace_cons_inv _ _)[σ2 [σ2' [? [?|[? Hsteps]]]]].
    + eexists σ2. split; [| by apply DemTraceUb].
      apply: (dem_has_trace_trans []) => //. by apply DemTraceUb.
    + have [? [??]]:= IH _ Hsteps => //.
      eexists. split => //.
      apply: (dem_has_trace_trans []) => //.
      by apply: DemTraceStep'.
Qed.

Lemma dem_has_trace_ub_app_inv {EV} κs (m : dem_module EV) σ1 σ2:
  σ1 ~{ m, κs ++ [Ub] }~>ₘ σ2 →
  ∃ σ3, σ1 ~{ m, κs }~>ₘ σ3 ∧ m.(dm_is_ub) σ3.
Proof.
  move => /dem_has_trace_app_inv[? [? /dem_has_trace_ub_inv [σ [??]]]].
  eexists σ. split; [ | done].
  apply: dem_has_trace_add_empty. by apply: dem_has_trace_trans.
Qed.

Program Definition dem_to_module {EV} (m : dem_module EV) := {|
  m_state := m.(dm_state);
  m_step σ e Pσ := (∃ σ', m.(dm_step) σ e σ' ∧ (∀ σ, Pσ σ ↔ σ = σ')) ∨ (m.(dm_is_ub) σ ∧ ¬ (∃ σ, Pσ σ));
|}.

Coercion dem_to_module : dem_module >-> module.

Lemma dem_has_trace_iff {EV} (m : dem_module EV) σ κs σ':
  σ ~{ m , κs }~>ₘ σ' ↔ σ ~{ m, κs }~> (σ' =.).
Proof.
  split.
  - elim.
    + move => ?. by constructor.
    + move => ? σ2 ??????.
      apply: (TraceStep (dem_to_module _) _ (σ2 =.)). { left. naive_solver. }
      naive_solver.
    + move => ????.
      apply: (TraceStep' _ _ (dem_to_module _) (λ _, False) _ _ None); [|done|naive_solver].
      right. naive_solver.
  - have : (∀ σ, eq σ' σ → eq σ' σ) by [].
    move: {1 3}(eq σ') => P HP Htrace.
    elim: Htrace HP.
    + move => σ2 ?? HP. rewrite (HP σ2) //. by constructor.
    + move => ????? [[?[??]]|[??]] ? IH ?.
      * apply: DemTraceStep; [done|]. apply: IH => //. naive_solver.
      * by apply: DemTraceUb.
Qed.

Lemma angelic_det_dem {EV} (m : dem_module EV):
  angelic_trace_det m.
Proof.
  move => ??? [[?[? HP]]|[??]].
  - right. eexists _. split => //. by apply HP. by move => ?? /HP -> ?.
  - by left.
Qed.

(*** properties of refines *)
Definition safe {EV} (m : mod_state EV) (P : list (event EV) → Prop) :=
  ∀ κs, m.(ms_state) ~{ m, κs }~> (λ _, True) → P κs.

Lemma refines_preserves_safe EV (mspec mimpl : mod_state EV) P:
  safe mspec P →
  mimpl ⊑ mspec →
  safe mimpl P.
Proof. move => Hs [Hr] κs Hκs. apply: Hs. by apply: Hr. Qed.

Global Instance refines_preorder EV : PreOrder (@refines EV).
Proof.
  constructor.
  - constructor => // κ Hi; naive_solver.
  - move => ??? [Hr1] [Hr2]. constructor => /=. naive_solver.
Qed.

(*** link *)
Record link_mediator EV1 EV2 EV3 := {
  lm_state : Type;
  lm_initial : lm_state;
  lm_step : lm_state → option EV1 → option EV2 → option EV3 → lm_state → Prop;
}.
Arguments lm_state {_ _ _}.
Arguments lm_initial {_ _ _}.
Arguments lm_step {_ _ _}.

Definition stateless_mediator {EV1 EV2 EV3} (R : option EV1 → option EV2 → option EV3 → Prop) : link_mediator EV1 EV2 EV3 := {|
  lm_state := unit;
  lm_initial := tt;
  lm_step _ e1 e2 e3 _:= R e1 e2 e3;
|}.

Inductive link_step {EV1 EV2 EV3} (m1 : module EV1) (m2 : module EV2) (M : link_mediator EV1 EV2 EV3) :
  m1.(m_state) * m2.(m_state) * M.(lm_state) → option EV3 → (m1.(m_state) * m2.(m_state) * M.(lm_state) → Prop) → Prop :=
| LinkStepL' σ1 σ2 e1 e' Pσ1' σm σm' (Pσ' : _ → Prop):
    m1.(m_step) σ1 e1 Pσ1' →
    (* TODO: is there a better way to formulate this? E.g. assume
    that there is no R None None Some in the theorem? *)
    (if e1 is Some es1 then M.(lm_step) σm e1 None e' σm' else e' = None ∧ σm' = σm) →
    (∀ σ', (Pσ1' σ'.1.1 ∧ σ'.1.2 = σ2 ∧ σ'.2 = σm') ↔ Pσ' σ') →
    link_step m1 m2 M (σ1, σ2, σm) e' Pσ'
| LinkStepR' σ1 σ2 e2 e' Pσ2' σm σm' (Pσ' : _ → Prop):
    m2.(m_step) σ2 e2 Pσ2' →
    (if e2 is Some es2 then M.(lm_step) σm None e2 e' σm' else e' = None ∧ σm' = σm) →
    (∀ σ', (σ'.1.1 = σ1 ∧ Pσ2' σ'.1.2 ∧ σ'.2 = σm') ↔ Pσ' σ') →
    link_step m1 m2 M (σ1, σ2, σm) e' Pσ'
| LinkStepBoth' σ1 σ2 e1 e2 e' Pσ1' Pσ2' σm σm' (Pσ' : _ → Prop):
    m1.(m_step) σ1 (Some e1) Pσ1' →
    m2.(m_step) σ2 (Some e2) Pσ2' →
    M.(lm_step) σm (Some e1) (Some e2) e' σm' →
    (∀ σ', (Pσ1' σ'.1.1 ∧ Pσ2' σ'.1.2 ∧ σ'.2 = σm') ↔ Pσ' σ') →
    link_step m1 m2 M (σ1, σ2, σm) e' Pσ'.

Lemma LinkStepL {EV1 EV2 EV3} (m1 : module EV1) (m2 : module EV2) (M : link_mediator EV1 EV2 EV3) σ1 σ2 e1 e' Pσ1' σm σm':
  m1.(m_step) σ1 e1 Pσ1' →
  (if e1 is Some es1 then M.(lm_step) σm e1 None e' σm' else e' = None ∧ σm' = σm) →
  link_step m1 m2 M (σ1, σ2, σm) e' (λ σ', Pσ1' σ'.1.1 ∧ σ'.1.2 = σ2 ∧ σ'.2 = σm' ).
Proof. move => ??. by apply: LinkStepL'. Qed.
Lemma LinkStepR {EV1 EV2 EV3} (m1 : module EV1) (m2 : module EV2) (M : link_mediator EV1 EV2 EV3) σ1 σ2 e2 e' Pσ2' σm σm':
  m2.(m_step) σ2 e2 Pσ2' →
  (if e2 is Some es2 then M.(lm_step) σm None e2 e' σm' else e' = None ∧ σm' = σm) →
  link_step m1 m2 M (σ1, σ2, σm) e' (λ σ', σ'.1.1 = σ1 ∧ Pσ2' σ'.1.2 ∧ σ'.2 = σm').
Proof. move => ??. by apply: LinkStepR'. Qed.
Lemma LinkStepBoth {EV1 EV2 EV3} (m1 : module EV1) (m2 : module EV2) (M : link_mediator EV1 EV2 EV3) σ1 σ2 e1 e2 e' Pσ1' Pσ2' σm σm':
  m1.(m_step) σ1 (Some e1) Pσ1' →
  m2.(m_step) σ2 (Some e2) Pσ2' →
  M.(lm_step) σm (Some e1) (Some e2) e' σm' →
  link_step m1 m2 M (σ1, σ2, σm) e' (λ σ', Pσ1' σ'.1.1 ∧ Pσ2' σ'.1.2 ∧ σ'.2 = σm').
Proof. move => ???. by apply: LinkStepBoth'. Qed.


Program Definition link {EV1 EV2 EV3} (m1 : module EV1) (m2 : module EV2) (M : link_mediator EV1 EV2 EV3) : module EV3 := {|
  m_state := m1.(m_state) * m2.(m_state) * M.(lm_state);
  m_step := (link_step m1 m2 M);
|}.

Lemma link_empty_steps_l {EV1 EV2 EV3} m1 m2 (M : link_mediator EV1 EV2 EV3) σ1 Pσ1' σ2 σm  :
  σ1 ~{ m1, [] }~> Pσ1' →
  (σ1, σ2, σm) ~{ link m1 m2 M, [] }~> (λ '(σ1', σ2', σm'), Pσ1' σ1' ∧ σ2' = σ2 ∧ σm = σm').
Proof.
  move Hκ: ([]) => κ Hsteps.
  elim: Hsteps Hκ.
  - move => ????. by apply: TraceEnd.
  - move => ??? [] //= ?????. apply: TraceStep'; [by apply: LinkStepL | done |].
    move => [[??]?] /= [?[??]]. naive_solver.
Qed.

Lemma link_empty_steps_r {EV1 EV2 EV3} m1 m2 (M : link_mediator EV1 EV2 EV3) σ1 Pσ2' σ2 σm :
  σ2 ~{ m2, [] }~> Pσ2' →
  (σ1, σ2, σm) ~{ link m1 m2 M, [] }~> (λ '(σ1', σ2', σm'), σ1' = σ1 ∧ Pσ2' σ2' ∧ σm = σm').
Proof.
  move Hκ: ([]) => κ Hsteps.
  elim: Hsteps Hκ.
  - move => ????. by apply: TraceEnd.
  - move => ??? [] //= ?????. apply: TraceStep'; [ by apply: LinkStepR | done | ].
    move => [[??]?] /= [?[??]]. naive_solver.
Qed.

(*
Inductive link_trace_related {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) : M.(lm_state) → list (event EV3) → (list (event EV1) → list (event EV2) → Prop) → Prop :=
| LinkTraceRelNil σm (Pκ : _ → _ → Prop):
    Pκ [] [] →
    link_trace_related M σm [] Pκ
| LinkTraceRelL (Pκ : _ → _ → Prop) Pκ' κ1 κ1' κs3 σm σm':
    M.(lm_step) σm (Some κ1) None κ1' σm' →
    (∀ κs1 κs2, Pκ κs1 κs2 → head κs1 = Some (Vis κ1) ∧ link_trace_related M σm' κs3 Pκ ∧ Pκ' (tail κs1) κs2) →
    link_trace_related M σm (option_list (Vis <$> κ1') ++ κs3) Pκ'.
(* | LinkTraceRelL κ1 κ1' κs1 κs2 κs3 σm σm': *)
(*     link_trace_related M σm' κs1 κs2 κs3 → *)
(*     M.(lm_step) σm (Some κ1) None κ1' σm' → *)
(*     link_trace_related M σm ([Vis κ1] ++ κs1) κs2 (option_list (Vis <$> κ1') ++ κs3) *)
(* | LinkTraceRelR κ2 κ2' κs1 κs2 κs3 σm σm': *)
(*     link_trace_related M σm' κs1 κs2 κs3 → *)
(*     M.(lm_step) σm None (Some κ2) κ2' σm' → *)
(*     link_trace_related M σm κs1 ([Vis κ2] ++ κs2) (option_list (Vis <$> κ2') ++ κs3) *)
(* | LinkTraceRelBoth κ1 κ2 κ3 κs1 κs2 κs3 σm σm': *)
(*     link_trace_related M σm' κs1 κs2 κs3 → *)
(*     M.(lm_step) σm (Some κ1) (Some κ2) κ3 σm' → *)
(*     link_trace_related M σm ([Vis κ1] ++ κs1) ([Vis κ2] ++ κs2) (option_list (Vis <$> κ3) ++ κs3) *)
(* . *)

Lemma link_trace_related_create {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) m1 m2 κs3 σ1 σ1':
  σ1 ~{ link m1 m2 M, κs3 }~> σ1' →
  link_trace_related M σ1.2 κs3 (λ κs1 κs2,
  σ1.1.1 ~{ m1, κs1 }~> (λ _, True) ∧
  σ1.1.2 ~{ m2, κs2 }~> (λ _, True)).
Proof. Admitted.
(*

  elim; clear.
  - move => σ Pσ ?. by econstructor; split; constructor.
  - move => σ1 Pσ2 Pσ3 κ κs Hstep Hsteps IH.
    inversion Hstep; clear Hstep; simplify_eq.
    + destruct e1; destruct_and?; simplify_eq/=.
      * apply: LinkTraceRelL; [done|].
        move => ???.

      have [?|[σ1[? Hκ1]]]:= HL1 _ _ _ ltac:(done).
      * eexists (option_list (Vis <$> e1) ++ [Ub]), [].
        split_and! => //;[ | | by apply: TraceEnd]; destruct e1; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //. by econstructor. }
        1: { econstructor. }
        all: apply: TraceStep'; [done..|] => ??; naive_solver.
      * have [|κs1 [κs2 [?[??]]]]:= IH (σ1, σ2, σm'); [ naive_solver|].
        eexists (option_list (Vis <$> e1) ++ κs1), κs2.
        split_and! => //; destruct e1; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
        all: apply: TraceStep'; [done..|] => ??.
        all: by apply: Hκ1; [..| done].
    + have [?|[σ[? Hκ2]]]:= HL2 _ _ _ ltac:(done).
      * eexists [], (option_list (Vis <$> e2) ++ [Ub]).
        split_and! => //;[ | by apply: TraceEnd |]; destruct e2; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //. by econstructor. }
        1: { econstructor. }
        all: apply: TraceStep'; [done..|] => ??; naive_solver.
      * have [|κs1 [κs2 [?[??]]]]:= IH (σ0, σ, σm'); [ naive_solver|].
        eexists κs1, (option_list (Vis <$> e2) ++ κs2).
        split_and! => //; destruct e2; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
        all: apply: TraceStep'; [done..|] => ??.
        all: by apply: Hκ2; [..| done].
    + have [?|[σ1[? Hκ1]]]:= HL1 _ _ _ ltac:(done). {
        eexists ([Vis e1; Ub]), [Vis e2].
        split_and! => //;[ | | apply: TraceStep' => // ??; apply: TraceEnd]; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //; by econstructor. }
        apply: TraceStep'; [done..|] => ??; naive_solver.
      }
      have [?|[σ[? Hκ2]]]:= HL2 _ _ _ ltac:(done). {
        eexists ([Vis e1]), [Vis e2; Ub].
        split_and! => //;[ | apply: TraceStep' => // ??; apply: TraceEnd |]; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //; by econstructor. }
        apply: TraceStep'; [done..|] => ??; naive_solver.
      }
      have [|κs1 [κs2 [?[??]]]]:= IH (σ1, σ, σm'); [ naive_solver|].
      eexists (Vis e1 :: κs1), (Vis e2 :: κs2).
      split_and! => //; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
      all: apply: TraceStep'; [done..|] => ??.
      all: try by apply: Hκ1; [..| done].
      all: try by apply: Hκ2; [..| done].
Qed.
 *)

Lemma link_trace_related_step {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) m1 m2 κs3 σ1 Pσ1' σ2 Pσ2' σm:
  link_trace_related M σm κs3 (λ κs1 κs2, σ1 ~{ m1, κs1 }~> Pσ1' ∧ σ2 ~{ m2, κs2 }~> Pσ2') →
  (σ1, σ2, σm) ~{ link m1 m2 M, κs3 }~> (λ '(σ1', σ2', σm''), Pσ1' σ1' ∧ Pσ2' σ2').
Proof.
  move => Hrel.
  elim: Hrel σ1 σ2. ; clear.
  - move => σm σ1 σ2 Hstep1 Hstep2. apply: (has_trace_trans [] []). { by apply: link_empty_steps_l. }
    move => [[??]?] [?[??]]. subst. apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?]?. apply: TraceEnd. naive_solver.
  - move => ????? /has_trace_ub_inv ? ?. apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?]. naive_solver.
  - move => ?????? /has_trace_ub_inv ?. apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?]. naive_solver.
  - move => κ1 κ1' κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= /(has_trace_cons_inv _ _)? ?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?] [[?[??]][??]]. subst. apply: TraceStep; [apply: LinkStepL; naive_solver|].
    move => [[??]?] /=[?[??]]. subst. apply: IH => //. naive_solver.
  - move => κ1 κ1' κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= ?/(has_trace_cons_inv _ _)?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?] [?[[?[??]]?]]. subst. apply: TraceStep; [apply: LinkStepR; naive_solver|].
    move => [[??]?] /=[?[??]]. subst. apply: IH => //. naive_solver.
  - move => κ1 κ2 κ3 κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= /(has_trace_cons_inv _ _)? /(has_trace_cons_inv _ _)?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?] [[?[??]][??]]. subst.
    apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?] [?[[?[??]]?]]. subst.
    apply: TraceStep; [ by apply: LinkStepBoth |].
    move => [[??]?] [?[??]]. subst.
    apply: IH => //; naive_solver.
Qed.

Lemma refines_horizontal {EV1 EV2 EV3} (m1 m2 m1' m2' : module _) σ1 σ2 σ1' σ2' (M : link_mediator EV1 EV2 EV3) :
  angelic_trace_det m1 →  angelic_trace_det m2 →
  MS m1 σ1 ⊑ MS m1' σ1' →
  MS m2 σ2 ⊑ MS m2' σ2' →
  MS (link m1 m2 M) (σ1, σ2, M.(lm_initial)) ⊑ MS (link m1' m2' M) (σ1', σ2', M.(lm_initial)).
Proof.
  move => ? ? [Hr1] [Hr2].
  constructor => κs /= /link_trace_related_create[//|//|?[?[?[??]]]].
  apply: has_trace_proper; [done..|].
  apply: link_trace_related_step => //.
  - by apply: Hr1.
  - by apply: Hr2.
Qed.
*)

(*
Inductive link_trace_related {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) : M.(lm_state) → list (event EV1) → list (event EV2) → list (event EV3) → Prop :=
| LinkTraceRelNil σm:
    link_trace_related M σm [] [] []
| LinkTraceRelUbL κs2 κs3 σm:
    link_trace_related M σm [Ub] κs2 κs3
| LinkTraceRelUbR κs1 κs3 σm:
    link_trace_related M σm κs1 [Ub] κs3
| LinkTraceRelL κ1 κ1' κs1 κs2 κs3 σm σm':
    link_trace_related M σm' κs1 κs2 κs3 →
    M.(lm_step) σm (Some κ1) None κ1' σm' →
    link_trace_related M σm ([Vis κ1] ++ κs1) κs2 (option_list (Vis <$> κ1') ++ κs3)
| LinkTraceRelR κ2 κ2' κs1 κs2 κs3 σm σm':
    link_trace_related M σm' κs1 κs2 κs3 →
    M.(lm_step) σm None (Some κ2) κ2' σm' →
    link_trace_related M σm κs1 ([Vis κ2] ++ κs2) (option_list (Vis <$> κ2') ++ κs3)
| LinkTraceRelBoth κ1 κ2 κ3 κs1 κs2 κs3 σm σm':
    link_trace_related M σm' κs1 κs2 κs3 →
    M.(lm_step) σm (Some κ1) (Some κ2) κ3 σm' →
    link_trace_related M σm ([Vis κ1] ++ κs1) ([Vis κ2] ++ κs2) (option_list (Vis <$> κ3) ++ κs3)
.

Lemma link_trace_related_create {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) m1 m2 κs3 σ1 σ1':
  angelic_trace_det m1 → angelic_trace_det m2 →
  σ1 ~{ link m1 m2 M, κs3 }~> σ1' →
  ∃ (Pκ : _ → _ → Prop), ∀ κs1 κs2, Pκ κs1 κs2 → link_trace_related M σ1.2 κs1 κs2 κs3 ∧
  σ1.1.1 ~{ m1, κs1 }~> (λ _, True) ∧
  σ1.1.2 ~{ m2, κs2 }~> (λ _, True).
Proof.
  move => HL1 HL2. elim; clear -HL1 HL2.
  - move => σ Pσ ?. eexists (λ κs1 κs2, κs1 = [] ∧ κs2 = []). move => ?? [-> ->]. by split_and!; constructor.
  - move => σ1 Pσ2 Pσ3 κ κs Hstep Hsteps IH.
    inversion Hstep; clear Hstep; simplify_eq.
    + eexists (λ κs1 κs2, ∃ σ2, Pσ2 σ2).
      move => ?? [??].

      have [?|[σ1[? Hκ1]]]:= HL1 _ _ _ ltac:(done).
      * eexists (option_list (Vis <$> e1) ++ [Ub]), [].
        split_and! => //;[ | | by apply: TraceEnd]; destruct e1; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //. by econstructor. }
        1: { econstructor. }
        all: apply: TraceStep'; [done..|] => ??; naive_solver.
      * have [|κs1 [κs2 [?[??]]]]:= IH (σ1, σ2, σm'); [ naive_solver|].
        eexists (option_list (Vis <$> e1) ++ κs1), κs2.
        split_and! => //; destruct e1; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
        all: apply: TraceStep'; [done..|] => ??.
        all: by apply: Hκ1; [..| done].
    + have [?|[σ[? Hκ2]]]:= HL2 _ _ _ ltac:(done).
      * eexists [], (option_list (Vis <$> e2) ++ [Ub]).
        split_and! => //;[ | by apply: TraceEnd |]; destruct e2; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //. by econstructor. }
        1: { econstructor. }
        all: apply: TraceStep'; [done..|] => ??; naive_solver.
      * have [|κs1 [κs2 [?[??]]]]:= IH (σ0, σ, σm'); [ naive_solver|].
        eexists κs1, (option_list (Vis <$> e2) ++ κs2).
        split_and! => //; destruct e2; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
        all: apply: TraceStep'; [done..|] => ??.
        all: by apply: Hκ2; [..| done].
    + have [?|[σ1[? Hκ1]]]:= HL1 _ _ _ ltac:(done). {
        eexists ([Vis e1; Ub]), [Vis e2].
        split_and! => //;[ | | apply: TraceStep' => // ??; apply: TraceEnd]; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //; by econstructor. }
        apply: TraceStep'; [done..|] => ??; naive_solver.
      }
      have [?|[σ[? Hκ2]]]:= HL2 _ _ _ ltac:(done). {
        eexists ([Vis e1]), [Vis e2; Ub].
        split_and! => //;[ | apply: TraceStep' => // ??; apply: TraceEnd |]; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //; by econstructor. }
        apply: TraceStep'; [done..|] => ??; naive_solver.
      }
      have [|κs1 [κs2 [?[??]]]]:= IH (σ1, σ, σm'); [ naive_solver|].
      eexists (Vis e1 :: κs1), (Vis e2 :: κs2).
      split_and! => //; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
      all: apply: TraceStep'; [done..|] => ??.
      all: try by apply: Hκ1; [..| done].
      all: try by apply: Hκ2; [..| done].
Qed.

Lemma link_trace_related_step {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) m1 m2 κs1 κs2 κs3 σ1 Pσ1' σ2 Pσ2' σm:
  link_trace_related M σm κs1 κs2 κs3 →
  σ1 ~{ m1, κs1 }~> Pσ1' →
  σ2 ~{ m2, κs2 }~> Pσ2' →
  (σ1, σ2, σm) ~{ link m1 m2 M, κs3 }~> (λ '(σ1', σ2', σm''), Pσ1' σ1' ∧ Pσ2' σ2').
Proof.
  move => Hrel.
  elim: Hrel σ1 σ2; clear.
  - move => σm σ1 σ2 Hstep1 Hstep2. apply: (has_trace_trans [] []). { by apply: link_empty_steps_l. }
    move => [[??]?] [?[??]]. subst. apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?]?. apply: TraceEnd. naive_solver.
  - move => ????? /has_trace_ub_inv ? ?. apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?]. naive_solver.
  - move => ?????? /has_trace_ub_inv ?. apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?]. naive_solver.
  - move => κ1 κ1' κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= /(has_trace_cons_inv _ _)? ?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?] [[?[??]][??]]. subst. apply: TraceStep; [apply: LinkStepL; naive_solver|].
    move => [[??]?] /=[?[??]]. subst. apply: IH => //. naive_solver.
  - move => κ1 κ1' κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= ?/(has_trace_cons_inv _ _)?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?] [?[[?[??]]?]]. subst. apply: TraceStep; [apply: LinkStepR; naive_solver|].
    move => [[??]?] /=[?[??]]. subst. apply: IH => //. naive_solver.
  - move => κ1 κ2 κ3 κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= /(has_trace_cons_inv _ _)? /(has_trace_cons_inv _ _)?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?] [[?[??]][??]]. subst.
    apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?] [?[[?[??]]?]]. subst.
    apply: TraceStep; [ by apply: LinkStepBoth |].
    move => [[??]?] [?[??]]. subst.
    apply: IH => //; naive_solver.
Qed.

Lemma refines_horizontal {EV1 EV2 EV3} (m1 m2 m1' m2' : module _) σ1 σ2 σ1' σ2' (M : link_mediator EV1 EV2 EV3) :
  angelic_trace_det m1 →  angelic_trace_det m2 →
  MS m1 σ1 ⊑ MS m1' σ1' →
  MS m2 σ2 ⊑ MS m2' σ2' →
  MS (link m1 m2 M) (σ1, σ2, M.(lm_initial)) ⊑ MS (link m1' m2' M) (σ1', σ2', M.(lm_initial)).
Proof.
  move => ? ? [Hr1] [Hr2].
  constructor => κs /= /link_trace_related_create[//|//|?[?[?[??]]]].
  apply: has_trace_proper; [done..|].
  apply: link_trace_related_step => //.
  - by apply: Hr1.
  - by apply: Hr2.
Qed.
*)
(*
Inductive link_trace_related {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) : M.(lm_state) → list (event EV1) → list (event EV2) → list (event EV3) → Prop :=
| LinkTraceRelNil σm:
    link_trace_related M σm [] [] []
| LinkTraceRelUbL κs2 κs3 σm:
    link_trace_related M σm [Ub] κs2 κs3
| LinkTraceRelUbR κs1 κs3 σm:
    link_trace_related M σm κs1 [Ub] κs3
| LinkTraceRelL κ1 κ1' κs1 κs2 κs3 σm σm':
    link_trace_related M σm' κs1 κs2 κs3 →
    M.(lm_step) σm (Some κ1) None κ1' σm' →
    link_trace_related M σm ([Vis κ1] ++ κs1) κs2 (option_list (Vis <$> κ1') ++ κs3)
| LinkTraceRelR κ2 κ2' κs1 κs2 κs3 σm σm':
    link_trace_related M σm' κs1 κs2 κs3 →
    M.(lm_step) σm None (Some κ2) κ2' σm' →
    link_trace_related M σm κs1 ([Vis κ2] ++ κs2) (option_list (Vis <$> κ2') ++ κs3)
| LinkTraceRelBoth κ1 κ2 κ3 κs1 κs2 κs3 σm σm':
    link_trace_related M σm' κs1 κs2 κs3 →
    M.(lm_step) σm (Some κ1) (Some κ2) κ3 σm' →
    link_trace_related M σm ([Vis κ1] ++ κs1) ([Vis κ2] ++ κs2) (option_list (Vis <$> κ3) ++ κs3)
.

Lemma link_trace_related_agree {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) m1 m2 κs1 κs2 κs3 σ1 σ2 σm Pσ Pσ1' κ:
  link_trace_related M σm κs1 κs2 κs3 →
  (σ1, σ2, σm) ~{ link m1 m2 M, κs3 }~> Pσ →
  m_step m1 σ1 κ Pσ1' →
  σ1 ~{ m1, κs1 }~> (λ _, True).
Proof.
Admitted.

Lemma link_trace_related_create {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) m1 m2 κs3 σ1 σ1':
  (* angelic_trace_det m1 → angelic_trace_det m2 → *)
  (∀ σ1 e Pσ1, m_step m1 σ1 e Pσ1 → LEM (∃ σ, Pσ1 σ)) →
  (∀ σ κs1, LEM (σ ~{ m1, κs1 }~> (λ _ : m_state m1, True))) →
  σ1 ~{ link m1 m2 M, κs3 }~> σ1' →
  ∃ κs1 κs2, link_trace_related M σ1.2 κs1 κs2 κs3 ∧
  σ1.1.1 ~{ m1, κs1 }~> (λ _, True) ∧
  σ1.1.2 ~{ m2, κs2 }~> (λ _, True).
Proof.
  move => HL1 HL2. elim; clear -HL1 HL2.
  - move => σ Pσ ?. eexists [], []. by split_and!; constructor.
  - move => σ1 Pσ2 Pσ3 κ κs Hstep Hsteps IH.
    inversion Hstep; clear Hstep; simplify_eq.
    + have [[σ?]|] := HL1 _ _ _ H.
      * have [|κs1[κs2[? [??]]]]:= IH (σ, σ2, σm'). naive_solver.
        eexists (option_list (Vis <$> e1) ++ κs1), κs2.
        split_and! => //; destruct e1; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
        all: apply: TraceStep'; [done..|] => σ1' ?.
        have ?:= Hsteps (σ1', σ2, σm') ltac:(naive_solver).
        have [//| Hσ1']:= HL2 σ1' κs1.
        exfalso.
        apply: link_trace_related_agree. done. done. done.

        all: by apply: Hκ1; [..| done].

      have [?|[σ1[? Hκ1]]]:= HL1 _ _ _ ltac:(done).
      * eexists (option_list (Vis <$> e1) ++ [Ub]), [].
        split_and! => //;[ | | by apply: TraceEnd]; destruct e1; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //. by econstructor. }
        1: { econstructor. }
        all: apply: TraceStep'; [done..|] => ??; naive_solver.
      * have [|κs1 [κs2 [?[??]]]]:= IH (σ1, σ2, σm'); [ naive_solver|].
        eexists (option_list (Vis <$> e1) ++ κs1), κs2.
        split_and! => //; destruct e1; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
        all: apply: TraceStep'; [done..|] => ??.
        all: by apply: Hκ1; [..| done].
    + have [?|[σ[? Hκ2]]]:= HL2 _ _ _ ltac:(done).
      * eexists [], (option_list (Vis <$> e2) ++ [Ub]).
        split_and! => //;[ | by apply: TraceEnd |]; destruct e2; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //. by econstructor. }
        1: { econstructor. }
        all: apply: TraceStep'; [done..|] => ??; naive_solver.
      * have [|κs1 [κs2 [?[??]]]]:= IH (σ0, σ, σm'); [ naive_solver|].
        eexists κs1, (option_list (Vis <$> e2) ++ κs2).
        split_and! => //; destruct e2; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
        all: apply: TraceStep'; [done..|] => ??.
        all: by apply: Hκ2; [..| done].
    + have [?|[σ1[? Hκ1]]]:= HL1 _ _ _ ltac:(done). {
        eexists ([Vis e1; Ub]), [Vis e2].
        split_and! => //;[ | | apply: TraceStep' => // ??; apply: TraceEnd]; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //; by econstructor. }
        apply: TraceStep'; [done..|] => ??; naive_solver.
      }
      have [?|[σ[? Hκ2]]]:= HL2 _ _ _ ltac:(done). {
        eexists ([Vis e1]), [Vis e2; Ub].
        split_and! => //;[ | apply: TraceStep' => // ??; apply: TraceEnd |]; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //; by econstructor. }
        apply: TraceStep'; [done..|] => ??; naive_solver.
      }
      have [|κs1 [κs2 [?[??]]]]:= IH (σ1, σ, σm'); [ naive_solver|].
      eexists (Vis e1 :: κs1), (Vis e2 :: κs2).
      split_and! => //; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
      all: apply: TraceStep'; [done..|] => ??.
      all: try by apply: Hκ1; [..| done].
      all: try by apply: Hκ2; [..| done].
Qed.

Lemma link_trace_related_step {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) m1 m2 κs1 κs2 κs3 σ1 Pσ1' σ2 Pσ2' σm:
  link_trace_related M σm κs1 κs2 κs3 →
  σ1 ~{ m1, κs1 }~> Pσ1' →
  σ2 ~{ m2, κs2 }~> Pσ2' →
  (σ1, σ2, σm) ~{ link m1 m2 M, κs3 }~> (λ '(σ1', σ2', σm''), Pσ1' σ1' ∧ Pσ2' σ2').
Proof.
  move => Hrel.
  elim: Hrel σ1 σ2; clear.
  - move => σm σ1 σ2 Hstep1 Hstep2. apply: (has_trace_trans [] []). { by apply: link_empty_steps_l. }
    move => [[??]?] [?[??]]. subst. apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?]?. apply: TraceEnd. naive_solver.
  - move => ????? /has_trace_ub_inv ? ?. apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?]. naive_solver.
  - move => ?????? /has_trace_ub_inv ?. apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?]. naive_solver.
  - move => κ1 κ1' κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= /(has_trace_cons_inv _ _)? ?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?] [[?[??]][??]]. subst. apply: TraceStep; [apply: LinkStepL; naive_solver|].
    move => [[??]?] /=[?[??]]. subst. apply: IH => //. naive_solver.
  - move => κ1 κ1' κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= ?/(has_trace_cons_inv _ _)?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?] [?[[?[??]]?]]. subst. apply: TraceStep; [apply: LinkStepR; naive_solver|].
    move => [[??]?] /=[?[??]]. subst. apply: IH => //. naive_solver.
  - move => κ1 κ2 κ3 κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= /(has_trace_cons_inv _ _)? /(has_trace_cons_inv _ _)?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?] [[?[??]][??]]. subst.
    apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?] [?[[?[??]]?]]. subst.
    apply: TraceStep; [ by apply: LinkStepBoth |].
    move => [[??]?] [?[??]]. subst.
    apply: IH => //; naive_solver.
Qed.

Lemma refines_horizontal {EV1 EV2 EV3} (m1 m2 m1' m2' : module _) σ1 σ2 σ1' σ2' (M : link_mediator EV1 EV2 EV3) :
  angelic_trace_det m1 →  angelic_trace_det m2 →
  MS m1 σ1 ⊑ MS m1' σ1' →
  MS m2 σ2 ⊑ MS m2' σ2' →
  MS (link m1 m2 M) (σ1, σ2, M.(lm_initial)) ⊑ MS (link m1' m2' M) (σ1', σ2', M.(lm_initial)).
Proof.
  move => ? ? [Hr1] [Hr2].
  constructor => κs /= /link_trace_related_create[//|//|?[?[?[??]]]].
  apply: has_trace_proper; [done..|].
  apply: link_trace_related_step => //.
  - by apply: Hr1.
  - by apply: Hr2.
Qed.
*)
Inductive link_trace_related {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) : M.(lm_state) → list (event EV1) → list (event EV2) → list (event EV3) → Prop :=
| LinkTraceRelNil σm:
    link_trace_related M σm [] [] []
| LinkTraceRelUbL κs2 κs3 σm:
    link_trace_related M σm [Ub] κs2 κs3
| LinkTraceRelUbR κs1 κs3 σm:
    link_trace_related M σm κs1 [Ub] κs3
| LinkTraceRelL κ1 κ1' κs1 κs2 κs3 σm σm':
    link_trace_related M σm' κs1 κs2 κs3 →
    M.(lm_step) σm (Some κ1) None κ1' σm' →
    link_trace_related M σm ([Vis κ1] ++ κs1) κs2 (option_list (Vis <$> κ1') ++ κs3)
| LinkTraceRelR κ2 κ2' κs1 κs2 κs3 σm σm':
    link_trace_related M σm' κs1 κs2 κs3 →
    M.(lm_step) σm None (Some κ2) κ2' σm' →
    link_trace_related M σm κs1 ([Vis κ2] ++ κs2) (option_list (Vis <$> κ2') ++ κs3)
| LinkTraceRelBoth κ1 κ2 κ3 κs1 κs2 κs3 σm σm':
    link_trace_related M σm' κs1 κs2 κs3 →
    M.(lm_step) σm (Some κ1) (Some κ2) κ3 σm' →
    link_trace_related M σm ([Vis κ1] ++ κs1) ([Vis κ2] ++ κs2) (option_list (Vis <$> κ3) ++ κs3)
.

Lemma link_trace_related_create {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) m1 m2 κs3 σ1 σ1':
  angelic_trace_det m1 → angelic_trace_det m2 →
  σ1 ~{ link m1 m2 M, κs3 }~> σ1' →
  ∃ κs1 κs2, link_trace_related M σ1.2 κs1 κs2 κs3 ∧
  σ1.1.1 ~{ m1, κs1 }~> (λ _, True) ∧
  σ1.1.2 ~{ m2, κs2 }~> (λ _, True).
Proof.
  move => HL1 HL2. elim; clear -HL1 HL2.
  - move => σ Pσ ?. eexists [], []. by split_and!; constructor.
  - move => σ1 Pσ2 Pσ3 κ κs Hstep Hsteps IH.
    inversion Hstep; clear Hstep; simplify_eq.
    + have [?|[σ1[? Hκ1]]]:= HL1 _ _ _ ltac:(done).
      * eexists (option_list (Vis <$> e1) ++ [Ub]), [].
        split_and! => //;[ | | by apply: TraceEnd]; destruct e1; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //. by econstructor. }
        1: { econstructor. }
        all: apply: TraceStep'; [done..|] => ??; naive_solver.
      * have [|κs1 [κs2 [?[??]]]]:= IH (σ1, σ2, σm'); [ naive_solver|].
        eexists (option_list (Vis <$> e1) ++ κs1), κs2.
        split_and! => //; destruct e1; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
        all: apply: TraceStep'; [done..|] => ??.
        all: by apply: Hκ1; [..| done].
    + have [?|[σ[? Hκ2]]]:= HL2 _ _ _ ltac:(done).
      * eexists [], (option_list (Vis <$> e2) ++ [Ub]).
        split_and! => //;[ | by apply: TraceEnd |]; destruct e2; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //. by econstructor. }
        1: { econstructor. }
        all: apply: TraceStep'; [done..|] => ??; naive_solver.
      * have [|κs1 [κs2 [?[??]]]]:= IH (σ0, σ, σm'); [ naive_solver|].
        eexists κs1, (option_list (Vis <$> e2) ++ κs2).
        split_and! => //; destruct e2; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
        all: apply: TraceStep'; [done..|] => ??.
        all: by apply: Hκ2; [..| done].
    + have [?|[σ1[? Hκ1]]]:= HL1 _ _ _ ltac:(done). {
        eexists ([Vis e1; Ub]), [Vis e2].
        split_and! => //;[ | | apply: TraceStep' => // ??; apply: TraceEnd]; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //; by econstructor. }
        apply: TraceStep'; [done..|] => ??; naive_solver.
      }
      have [?|[σ[? Hκ2]]]:= HL2 _ _ _ ltac:(done). {
        eexists ([Vis e1]), [Vis e2; Ub].
        split_and! => //;[ | apply: TraceStep' => // ??; apply: TraceEnd |]; destruct_and?; simplify_eq/= => //; rewrite ?right_id //.
        1: { econstructor => //; by econstructor. }
        apply: TraceStep'; [done..|] => ??; naive_solver.
      }
      have [|κs1 [κs2 [?[??]]]]:= IH (σ1, σ, σm'); [ naive_solver|].
      eexists (Vis e1 :: κs1), (Vis e2 :: κs2).
      split_and! => //; destruct_and?; simplify_eq/= => //; rewrite ?right_id //. by econstructor.
      all: apply: TraceStep'; [done..|] => ??.
      all: try by apply: Hκ1; [..| done].
      all: try by apply: Hκ2; [..| done].
Qed.

Lemma link_trace_related_step {EV1 EV2 EV3} (M : link_mediator EV1 EV2 EV3) m1 m2 κs1 κs2 κs3 σ1 Pσ1' σ2 Pσ2' σm:
  link_trace_related M σm κs1 κs2 κs3 →
  σ1 ~{ m1, κs1 }~> Pσ1' →
  σ2 ~{ m2, κs2 }~> Pσ2' →
  (σ1, σ2, σm) ~{ link m1 m2 M, κs3 }~> (λ '(σ1', σ2', σm''), Pσ1' σ1' ∧ Pσ2' σ2').
Proof.
  move => Hrel.
  elim: Hrel σ1 σ2; clear.
  - move => σm σ1 σ2 Hstep1 Hstep2. apply: (has_trace_trans [] []). { by apply: link_empty_steps_l. }
    move => [[??]?] [?[??]]. subst. apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?]?. apply: TraceEnd. naive_solver.
  - move => ????? /has_trace_ub_inv ? ?. apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?]. naive_solver.
  - move => ?????? /has_trace_ub_inv ?. apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?]. naive_solver.
  - move => κ1 κ1' κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= /(has_trace_cons_inv _ _)? ?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?] [[?[??]][??]]. subst. apply: TraceStep; [apply: LinkStepL; naive_solver|].
    move => [[??]?] /=[?[??]]. subst. apply: IH => //. naive_solver.
  - move => κ1 κ1' κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= ?/(has_trace_cons_inv _ _)?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?] [?[[?[??]]?]]. subst. apply: TraceStep; [apply: LinkStepR; naive_solver|].
    move => [[??]?] /=[?[??]]. subst. apply: IH => //. naive_solver.
  - move => κ1 κ2 κ3 κs1 κs2 κs3 ?? ? IH HR σ1 σ2 /= /(has_trace_cons_inv _ _)? /(has_trace_cons_inv _ _)?.
    apply: (has_trace_trans []). { by apply: link_empty_steps_l. }
    move => [[??]?] [[?[??]][??]]. subst.
    apply: (has_trace_trans []). { by apply: link_empty_steps_r. }
    move => [[??]?] [?[[?[??]]?]]. subst.
    apply: TraceStep; [ by apply: LinkStepBoth |].
    move => [[??]?] [?[??]]. subst.
    apply: IH => //; naive_solver.
Qed.

Lemma refines_horizontal {EV1 EV2 EV3} (m1 m2 m1' m2' : module _) σ1 σ2 σ1' σ2' (M : link_mediator EV1 EV2 EV3) :
  angelic_trace_det m1 →  angelic_trace_det m2 →
  MS m1 σ1 ⊑ MS m1' σ1' →
  MS m2 σ2 ⊑ MS m2' σ2' →
  MS (link m1 m2 M) (σ1, σ2, M.(lm_initial)) ⊑ MS (link m1' m2' M) (σ1', σ2', M.(lm_initial)).
Proof.
  move => ? ? [Hr1] [Hr2].
  constructor => κs /= /link_trace_related_create[//|//|?[?[?[??]]]].
  apply: has_trace_proper; [done..|].
  apply: link_trace_related_step => //.
  - by apply: Hr1.
  - by apply: Hr2.
Qed.
(*** has_non_ub_trace *)
Inductive has_non_ub_trace {EV} (m : dem_module EV) : m.(dm_state) → list EV → m.(dm_state) → Prop :=
| NUBTraceEnd σ:
    has_non_ub_trace m σ [] σ
| NUBTraceStep σ1 σ2 σ3 κ κs:
    m.(dm_step) σ1 κ σ2 →
    has_non_ub_trace m σ2 κs σ3 →
    has_non_ub_trace m σ1 (option_list κ ++ κs) σ3
.
Notation " σ '~{' m , κ '}~>ₙ' σ' " := (has_non_ub_trace m σ κ σ') (at level 40).
Notation " σ '~{' m , κ '}~>ₙ' - " := (∃ σ', has_non_ub_trace m σ κ σ') (at level 40).

Lemma NUBTraceStepNone {EV} κs (m : dem_module EV) σ2 σ1 σ3 :
  m.(dm_step) σ1 None σ2 →
  σ2 ~{ m, κs }~>ₙ σ3 →
  σ1 ~{ m, κs }~>ₙ σ3.
Proof. move => ??. by apply: (NUBTraceStep _ _ _ _ None). Qed.

Lemma NUBTraceStepSome {EV} κs (m : dem_module EV) σ2 σ1 σ3 κ :
  m.(dm_step) σ1 (Some κ) σ2 →
  σ2 ~{ m, κs }~>ₙ σ3 →
  σ1 ~{ m, κ :: κs }~>ₙ σ3.
Proof. move => ??. by apply: (NUBTraceStep _ _ _ _ (Some _)). Qed.

Lemma has_non_ub_trace_trans {EV} κs1 κs2 (m : dem_module EV) σ1 σ2 σ3 :
  σ1 ~{ m, κs1 }~>ₙ σ2 →
  σ2 ~{ m, κs2 }~>ₙ σ3 →
  σ1 ~{ m, κs1 ++ κs2 }~>ₙ σ3.
Proof.
  elim => //.
  move => ?????????. rewrite -app_assoc. econstructor; eauto.
Qed.

Lemma has_non_ub_trace_add_empty {EV} κs1 (m : dem_module EV) σ1 σ2 :
  σ1 ~{ m, κs1 ++ [] }~>ₙ σ2 →
  σ1 ~{ m, κs1 }~>ₙ σ2.
Proof. by rewrite -{2}[κs1](right_id_L [] (++)). Qed.

Lemma has_trace_to_non_ub_trace EV (m : dem_module EV) σ1 κs σ2:
  σ1 ~{ m, κs }~>ₘ σ2 →
  ∃ κs' σ2', Vis <$> κs' `prefix_of` κs ∧ σ1 ~{ m, κs' }~>ₙ σ2' ∧
             ((Vis <$> κs' = κs ∧ σ2' = σ2) ∨ m.(dm_is_ub) σ2').
Proof.
  elim.
  - move => ?. eexists [], _. naive_solver constructor.
  - move => ??? κ ??? [κs' [σ2' [?[??]]]]. eexists (option_list κ ++ κs'), σ2'.
    split_and! => //.
    + destruct κ => //. by apply: prefix_cons.
    + by econstructor.
    + destruct κ; naive_solver.
  - move => ????. eexists [], _. split_and! => //=.
    + by apply prefix_nil.
    + by constructor.
    + by right.
Qed.

(*** has_no_behavior *)
Definition has_no_behavior {EV} (m : module EV) (σ : m.(m_state)) :=
  ∀ σ' κs, σ ~{ m, κs }~> σ' → κs = [].

Lemma no_behavior_step {EV} (m : module EV) σ:
  (∀ e Pσ', m.(m_step) σ e Pσ' → e = None ∧ ∃ σ', Pσ' σ' ∧ has_no_behavior m σ') →
  has_no_behavior m σ.
Proof.
  move => Hstep ?? Htrace. inversion Htrace; simplify_eq/= => //.
  have [-> [? [? Hnext]]] := Hstep _ _ H => /=. apply: Hnext. naive_solver.
Qed.

(*** state_set *)
Definition state_set_refines {EV} (mimpl mspec : module EV) (σi : mimpl.(m_state)) (σs : propset mspec.(m_state)) : Prop :=
  ∀ κs, σi ~{ mimpl, κs }~> (λ _, True) → ∃ σs1, σs1 ∈ σs ∧ σs1 ~{ mspec, κs }~> (λ _, True).

Lemma inv_set_implies_refines {EV} (m1 m2 : mod_state EV) (inv : m1.(m_state) → propset m2.(m_state) → Prop):
  inv m1.(ms_state) {[ m2.(ms_state) ]} →
  (∀ σi σs, inv σi σs → ∃ σ, σ ∈ σs) →
  (* (∀ σi σs, inv σi σs → m1.(m_is_ub) σi → ∃ σs1, σs1 ∈ σs ∧ σs1 ~{ m2, [Ub] }~> (λ _, True)) → *)
  (* (∀ σi1 σs1 σi2 e, inv σi1 σs1 → m1.(m_step) σi1 e σi2 → *)
      (* ∃ σs2, inv σi2 σs2 ∧ σs2 ⊆ {[ σ2 | ∃ σ1, σ1 ∈ σs1 ∧ σ1 ~{ m2, option_list (Vis <$> e) }~> σ2 ]}) → *)
  (∀ σi1 σs1 Pσi2 e, inv σi1 σs1 → m1.(m_step) σi1 e Pσi2 → ∃ σs2, ∀ σi2, inv σi2 σs2 ∧ (Pσi2 σi2 →
      ∃ σ1, σ1 ∈ σs1 ∧ σ1 ~{ m2, option_list (Vis <$> e) }~> (λ x, x ∈ σs2))) →
  m1 ⊑ m2.
Proof.
  move => Hinvinit Hinvnonempty Hinvstep.
  constructor => // κs.
  move: m1.(ms_state) Hinvinit => σi1 Hinv Hsteps.
  have : (∃ σs1, σs1 ∈ ({[ms_state m2]} : propset _) ∧ σs1 ~{ m2, κs }~> (λ _, True)); last set_solver.
  move: {[ m2.(ms_state) ]} Hinv => σs1 Hinv.
  elim: Hsteps σs1 Hinv => {σi1 κs}.
  - move => ???? /Hinvnonempty [??]. eexists _. split => //. by apply: TraceEnd.
  - move => σi1 σi2 σi3 κ κs Hstep Hsteps IH σs1 Hinv.
    have := Hinvstep _ _ _ _ Hinv Hstep.
    (* TODO: continue here. The lemma statement is probably wrong *)

    have [σs2 [Hinv2 Hsub]]:= Hinvstep _ _ _ _ Hinv Hstep.
    have [σs3 [σs4 [Hin ?]]]:= IH _ Hinv2.
    have [σ1 [??]]:= Hsub _ Hin.
    eexists _, _. split => //. by apply: has_trace_trans.
  - move => ??? /Hinvsafe Hs σs Hinv.
    have [? [? [? /has_trace_ub_inv[σs2[??]]]]]:= Hs _ Hinv.
    eexists _, _. split => //. apply: (has_trace_trans []); [ done |]. by apply: TraceUbRefl.
Qed.
  move => Hinvinit Hinvnonempty Hinvsafe Hinvstep.
  constructor => // κs [σi2].
  move: m1.(ms_state) Hinvinit => σi1 Hinv Hsteps.
  have : (∃ σs1 σs2, σs1 ∈ ({[ms_state m2]} : propset _) ∧ σs1 ~{ m2, κs }~> σs2); last set_solver.
  move: {[ m2.(ms_state) ]} Hinv => σs1 Hinv.
  elim: Hsteps σs1 Hinv => {σi1 σi2 κs}.
  - move => ? ? /Hinvnonempty [??].  eexists _, _. split => //. by apply: TraceEnd.
  - move => σi1 σi2 σi3 κ κs Hstep Hsteps IH σs1 Hinv.
    have [σs2 [Hinv2 Hsub]]:= Hinvstep _ _ _ _ Hinv Hstep.
    have [σs3 [σs4 [Hin ?]]]:= IH _ Hinv2.
    have [σ1 [??]]:= Hsub _ Hin.
    eexists _, _. split => //. by apply: has_trace_trans.
  - move => ??? /Hinvsafe Hs σs Hinv.
    have [? [? [? /has_trace_ub_inv[σs2[??]]]]]:= Hs _ Hinv.
    eexists _, _. split => //. apply: (has_trace_trans []); [ done |]. by apply: TraceUbRefl.
Qed.

Lemma state_set_refines_initial {EV} (m1 m2 : mod_state EV):
  m1 ⊑ m2 →
  state_set_refines m1 m2 (ms_state m1) {[ms_state m2]}.
Proof. move => Hr ?? /(refines_explicit _ m2)[//|??]. naive_solver. Qed.

Lemma state_set_refines_step {EV} (m1 m2 : module EV) σi1 σs1 σi2 e:
  state_set_refines m1 m2 σi1 σs1 →
  m1.(m_step) σi1 e σi2 →
  state_set_refines m1 m2 σi2 {[ σ2 | ∃ σ1, σ1 ∈ σs1 ∧ σ1 ~{ m2, option_list (Vis <$> e) }~> σ2 ]}.
Proof.
  move => Hinv Hstep κs σi3 Hκs.
  have [|? [? [? /has_trace_app_inv[?[??]]]]]:= Hinv (option_list (Vis <$> e) ++ κs) σi3.
  { by apply: TraceStep. }
  set_solver.
Qed.

Lemma state_set_refines_step_None {EV} (m1 m2 : module EV) σi1 σs1 σi2:
  state_set_refines m1 m2 σi1 σs1 →
  m1.(m_step) σi1 None σi2 →
  state_set_refines m1 m2 σi2 σs1.
Proof.
  move => Hinv Hstep κs σi3 Hκs.
  have [|? [? [? ?]]]:= Hinv κs σi3.
  { by apply: TraceStepNone. }
  set_solver.
Qed.

Lemma state_set_refines_non_empty {EV} (m1 m2 : module EV) σi σs:
  state_set_refines m1 m2 σi σs → ∃ σ, σ ∈ σs.
Proof.
  move => Hs.
  have [|?[?[??]]]:= Hs [] σi. by apply: TraceEnd.
  naive_solver.
Qed.

Lemma state_set_refines_ub {EV} (m1 m2 : module EV) σi σs:
  state_set_refines m1 m2 σi σs →
  m1.(m_is_ub) σi →
  ∃ σ, σ ∈ σs ∧ σ ~{ m2, [Ub] }~> -.
Proof. move => Hs Hub. apply: Hs. by apply: TraceUbRefl. Qed.

Lemma refines_implies_inv_set {EV} (m1 m2 : mod_state EV):
  m1 ⊑ m2 →
  ∃ (inv : m1.(m_state) → propset m2.(m_state) → Prop),
  inv m1.(ms_state) {[ m2.(ms_state) ]} ∧
  (∀ σi σs, inv σi σs → ∃ σ, σ ∈ σs) ∧
  (∀ σi σs, inv σi σs → m1.(m_is_ub) σi → ∃ σs1, σs1 ∈ σs ∧ σs1 ~{ m2, [Ub] }~> -) ∧
  (∀ σi1 σs1 σi2 e, inv σi1 σs1 → m1.(m_step) σi1 e σi2 →
      ∃ σs2, inv σi2 σs2 ∧ σs2 ⊆ {[ σ2 | ∃ σ1, σ1 ∈ σs1 ∧ σ1 ~{ m2, option_list (Vis <$> e) }~> σ2 ]}).
Proof.
  move => Href.
  eexists (state_set_refines m1 m2).
  split_and!.
  - by apply: state_set_refines_initial.
  - by apply: state_set_refines_non_empty.
  - move => σi σs Hinv Hub. by apply: state_set_refines_ub.
  - move => σi1 σs1 σi2 e Hinv Hstep.
    eexists _. split_and!; last reflexivity.
    by apply: state_set_refines_step.
Qed.

(*** wp': equivalent definition of refines *)
Inductive wp' {EV} (m1 : module EV) (m2 : mod_state EV) : nat → m1.(m_state) -> list (event EV) -> Prop :=
| Wp_step' σi1 κs n:
     (∃ σs2, m2.(ms_state) ~{ m2, κs }~> σs2 ∧ m2.(m_is_ub) σs2) ∨
       ¬ m1.(m_is_ub) σi1 ∧
       (∀ σi2 κ n', n = S n' → m1.(m_step) σi1 κ σi2 ->
         ∃ σs2, m2.(ms_state) ~{ m2, κs ++ option_list (Vis <$> κ) }~> σs2 ∧
               wp' m1 m2 n' σi2 (κs ++ option_list (Vis <$> κ))) ->
    wp' m1 m2 n σi1 κs
.

Lemma wp'_weaken {EV} (m1 : module EV) m2 κs σ n n':
  n' ≤ n →
  wp' m1 m2 n σ κs →
  wp' m1 m2 n' σ κs.
Proof.
  elim: n' n σ κs.
  - move => ???? Hwp. constructor.
    inversion Hwp as [??? Hwp']; simplify_eq. have [|[? _]]:= Hwp'. naive_solver.
    right. split; [ done | lia].
  - move => n' IH [|n] σ κs ? Hwp. lia.
    inversion Hwp as [??? Hwp']; simplify_eq.
    constructor.
    have [|[? {}Hwp']]:= Hwp'. naive_solver.
    right. split => // σi2 κ n'' [?] ?. subst.
    have [//|? [? ?]]:= Hwp' σi2 κ _ ltac:(done).
    eexists. split => //. apply: IH; [|done]. lia.
Qed.

Lemma forall_to_ex A B (P : A → B → Prop) (Q : B → Prop):
 (∃ n : A, ∀ y : B, P n y → Q y) -> ∀ y : B, ((∀ n : A, P n y) → Q y).
Proof. naive_solver. Qed.

Lemma wp'_implies_refines {EV} (m1 m2 : mod_state EV):
  (∀ n, wp' m1 m2 n m1.(ms_state) []) →
  m1 ⊑ m2.
Proof.
  move => Hwp.
  constructor => κs [σi].
  move: m1.(ms_state) Hwp => σi1.
  have : (has_trace m2 m2.(ms_state) [] m2.(ms_state)). { by apply: TraceEnd. }
  move: {2}m2.(ms_state) => σs1.
  have : κs = [] ++ κs by [].
  move: ([]) => κstart. move: {2 3}(κs) => κend.
  move => Hκ Hs Hwp Hsteps.
  move: κstart Hwp σs1 Hs Hκ. apply: forall_to_ex.
  elim: Hsteps => {σi1 κend σi}.
  - move => σi1. exists 0 => κstart Hwp σs Hs Hκ.
    rewrite right_id in Hκ; subst. naive_solver.
  - move => σi1 σi2 σi3 κ κend Hstep Hsteps [n IH]. exists (S n) => κstart Hwp σs1 Hs Hκs.
    inversion_clear Hwp as [??? Hwp2]; subst.
    case: Hwp2 => [[σs [Hub1 Hub2]]|[? {} Hwp]]. {
      eexists σs. apply: has_trace_trans => //. by apply: TraceUb.
    }
    have [|σs2 [Hsteps2 {}Hwp]]:= (Hwp _ _ n _ Hstep) => //.
    have [|??]:= (IH _ Hwp _ Hsteps2) => //. by rewrite assoc.
    by eexists.
  - move => σ1 ???. exists 0 => ? Hwp ???.
    inversion_clear Hwp as [??? Hwp2]; subst.
    case: Hwp2 => [[σs [Hub1 Hub2]]|[? //]].
    eexists σs. apply: has_trace_trans => //. by apply: TraceUb.
Qed.

Lemma refines_implies_wp' {EV} (m1 m2 : mod_state EV):
  (∀ σ, LEM (m1.(m_is_ub) σ)) →
  m1 ⊑ m2 →
  (∀ n, wp' m1 m2 n m1.(ms_state) []).
Proof.
  move => Hdec Hr n.
  have : (has_trace m1 m1.(ms_state) [] m1.(ms_state)). { by apply: TraceEnd. }
  move: {2 3}(m1.(ms_state)) => σi.
  move: ([]) => κstart.
  elim/lt_wf_ind: n κstart σi.
  move => n IH κstart σi Hstepi.
  constructor.
  have [??]:= (refines_explicit _ _ _ _ Hr Hstepi).
  have [?|?] := Hdec σi. {
    left.
    have /(refines_explicit _ _ _ _ Hr)[? /has_trace_ub_app_inv ? //]: has_trace m1 (ms_state m1) (κstart ++ [Ub]) σi.
    apply: has_trace_trans => //. by apply: TraceUb.
  }
  right. split => // σi2 κ n' ? Hstep; subst.
  have Hs1' : has_trace m1 (ms_state m1) (κstart ++ option_list (Vis <$> κ)) σi2. {
    apply: has_trace_trans => //.
    rewrite -(right_id_L [] (++) (option_list _)).
    apply: TraceStep => //. by apply: TraceEnd.
  }
  move: (Hs1') => /(refines_explicit _ _ _ _ Hr)[??].
  eexists _. split => //.
  apply: IH => //. lia.
Qed.

(*** Proving refinement *)
Lemma inv_implies_refines {EV} (m1 m2 : mod_state EV) (inv : m1.(m_state) → m2.(m_state) → Prop):
  inv m1.(ms_state) m2.(ms_state) →
  (∀ σi σs, inv σi σs → ¬ m1.(m_is_ub) σi) →
  (∀ σi1 σs1 σi2 e,
      inv σi1 σs1 → m1.(m_step) σi1 e σi2 →
      ∃ σs2, σs1 ~{ m2, option_list (Vis <$> e) ++ [Ub] }~> σs2 ∨ (inv σi2 σs2 ∧ σs1 ~{ m2, option_list (Vis <$> e) }~> σs2)) →
  m1 ⊑ m2.
Proof.
  move => Hinvinit Hinvsafe Hinvstep.
  constructor => // κs [σi2]. move: m1.(ms_state) m2.(ms_state) Hinvinit => σi1 σs1 Hinv Hsteps.
  elim: Hsteps σs1 Hinv => {σi1 σi2 κs}.
  - by eauto using TraceEnd.
  - move => σi1 σi2 σi3 κ κs Hstep Hsteps IH σs1 Hinv.
    case: (Hinvstep _ _ _ _ Hinv Hstep) => σs2 [/has_trace_app_inv [? [? /has_trace_ub_inv [σub [? ?]]]]|[Hinv2 ?]]. {
      eexists σs2. apply: has_trace_trans => //. apply: (has_trace_trans []) => //. by apply: TraceUb.
    }
    case: (IH _ Hinv2) => ? ?.
    eexists. by apply: has_trace_trans.
  - move => ??? /Hinvsafe ? σs ?. exists σs. naive_solver.
Qed.

Lemma inv_implies_refines' {EV} (m1 m2 : mod_state EV) (inv : m1.(m_state) → m2.(m_state) → Prop):
  inv m1.(ms_state) m2.(ms_state) →
  (∀ σi σs, inv σi σs → m1.(m_is_ub) σi → ∃ σs2, σs ~{ m2, [Ub] }~> σs2) →
  (∀ σi1 σs1 σi2 e, inv σi1 σs1 → m1.(m_step) σi1 e σi2 →
      (m1.(m_is_ub) σi1 ∨ m2.(m_is_ub) σs1) ∨
      ∃ σs2, (inv σi2 σs2 ∨ has_no_behavior m1 σi2) ∧ σs1 ~{ m2, option_list (Vis <$> e) }~> σs2) →
  m1 ⊑ m2.
Proof.
  move => Hinvinit Hinvsafe Hinvstep.
  constructor => // κs [σi2].
  move: m1.(ms_state) m2.(ms_state) Hinvinit => σi1 σs1 Hinv Hsteps.
  elim: Hsteps σs1 Hinv => {σi1 σi2 κs}.
  - by eauto using TraceEnd.
  - move => σi1 σi2 σi3 κ κs Hstep Hsteps IH σs1 Hinv.
    case: (Hinvstep _ _ _ _ Hinv Hstep) => [|[σs2 [Hinv2 ?]]]. {
      case => Hub; [|eexists _; by apply: TraceUbRefl].
      have [? /has_trace_ub_inv[σs2[??]]]:= Hinvsafe _ _ Hinv Hub.
      eexists σs2. apply: (has_trace_trans []); [ done |]. by apply: TraceUb.
    }
    case: Hinv2 => Hinv2. 2: {
      eexists _. apply: has_trace_trans => //.
      have -> := Hinv2 _ _ Hsteps.
        by apply: TraceEnd.
    }
    case: (IH _ Hinv2) => ? ?.
    eexists. by apply: has_trace_trans.
  - move => ??? /Hinvsafe Hs σs Hinv. have [? /has_trace_ub_inv[σs2[??]]]:= Hs _ Hinv.
    eexists σs2. apply: (has_trace_trans []); [ done |]. by apply: TraceUb.
Qed.

(* This does not seem nice to work work. *)
Lemma inv_implies_refines_equiv {EV} (m1 m2 : mod_state EV) (inv : m1.(m_state) → m2.(m_state) → Prop):
  inv m1.(ms_state) m2.(ms_state) →
  (∀ σi σs, inv σi σs → m1.(m_is_ub) σi → ∃ σs2, σs ~{ m2, [Ub] }~> σs2) →
  (∀ σi σs, inv σs σi → m2.(m_is_ub) σi → ∃ σs2, σs ~{ m1, [Ub] }~> σs2) →
  (∀ σi1 σs1 σi2 e, inv σi1 σs1 → m1.(m_step) σi1 e σi2 →
      (m1.(m_is_ub) σi1 ∨ m2.(m_is_ub) σs1) ∨
      ∃ σs2, (inv σi2 σs2 ∨ has_no_behavior m1 σi2) ∧ σs1 ~{ m2, option_list (Vis <$> e) }~> σs2) →
  (∀ σi1 σs1 σs2 e, inv σi1 σs1 → m2.(m_step) σs1 e σs2 →
      (m1.(m_is_ub) σi1 ∨ m2.(m_is_ub) σs1) ∨
      ∃ σi2, (inv σi2 σs2 ∨ has_no_behavior m2 σs2) ∧ σi1 ~{ m1, option_list (Vis <$> e) }~> σi2) →
  refines_equiv m1 m2.
Proof.
  move => Hinvinit Hinvsafe1 Hinvsafe2 Hinvstep1 Hinvstep2.
  split; [ apply: inv_implies_refines' => //; naive_solver |].
  apply: (inv_implies_refines' _ _ (flip inv)) => //=; naive_solver.
Qed.

(* This does not seem nice to work work. *)
(* Lemma link_merge_calls {EV1 EV2 EV3} (m1 : module EV1) (m2 : module EV2) (m3 : module EV3) (inv : m1.(m_state) → m2.(m_state) → m3.(m_state) → Prop) R : *)
(*   let R' e1 e2 e3 := if (e1, e2) is (None, None) then e3 = None else R e1 e2 e3 in *)
(*   inv m1.(m_initial) m2.(m_initial) m3.(m_initial) → *)
(*   (∀ σ1 σ2 σ3, inv σ1 σ2 σ3 → m3.(m_is_ub) σ3 ↔ (m1.(m_is_ub) σ1 ∨ m2.(m_is_ub) σ2)) → *)
(*   (∀ σ1 σ2 σ3, inv σ1 σ2 σ3 → ∀ e σ32, m_step m3 σ3 e σ32 → ∃ σ12 σ22, link_step m1 m2 R (σ1, σ2) e (σ12, σ22) ∧ inv σ12 σ22 σ32) → *)
(*   (∀ σ1 σ2 σ3, inv σ1 σ2 σ3 → ∀ e σ12 e', m_step m1 σ1 e σ12 → R' e None e' → ∃ σ32, m3.(m_step) σ3 e' σ32 ∧ inv σ12 σ2 σ32) → *)
(*   (∀ σ1 σ2 σ3, inv σ1 σ2 σ3 → ∀ e σ22 e', m_step m2 σ2 e σ22 → R' None e e' → ∃ σ32, m3.(m_step) σ3 e' σ32 ∧ inv σ1 σ22 σ32) → *)
(*   (∀ σ1 σ2 σ3, inv σ1 σ2 σ3 → ∀ e1 e2 σ12 σ22 e', m_step m1 σ1 (Some e1) σ12 → m_step m2 σ2 (Some e2) σ22 → R (Some e1) (Some e2) e' → ∃ σ32, m3.(m_step) σ3 e' σ32 ∧ inv σ12 σ22 σ32) → *)
(*   refines_equiv (link m1 m2 R) m3. *)
(* Proof. *)
(*   move => R' Hinit Hub Hmstep3 Hmstep1 Hmstep2 Hmstepboth. *)
(*   apply: (inv_implies_refines_equiv (link m1 m2 R) m3 (λ '(σ1, σ2) σ3, inv σ1 σ2 σ3)). *)
(*   - done. *)
(*   - move => [??] ?. naive_solver. *)
(*   - move => [σ11 σ21] σ31 [σ12 σ22] e Hinv Hstep. inversion Hstep; simplify_eq/=. *)
(*     + revert select (m_step _ _ _ _) => /(Hmstep1 _ _ _ Hinv) Hm3. *)
(*       destruct e1; simplify_eq; move: (Hm3 _ ltac:(done)) => [σ32 [? ?]]. *)
(*       all: eexists σ32; split => //; apply: has_trace_add_empty; apply: TraceStep => //; by apply: TraceEnd. *)
(*     + revert select (m_step _ _ _ _) => /(Hmstep2 _ _ _ Hinv) Hm3. *)
(*       destruct e2; simplify_eq; move: (Hm3 _ ltac:(done)) => [σ32 [? ?]]. *)
(*       all: eexists σ32; split => //; apply: has_trace_add_empty; apply: TraceStep => //; by apply: TraceEnd. *)
(*     + revert select (m_step _ _ _ _) => /(Hmstepboth _ _ _ Hinv) Hm3. *)
(*       revert select (m_step _ _ _ _) => /Hm3 {}Hm3. *)
(*       revert select (R _ _ _) => /Hm3 [σ32 [? ?]]. *)
(*       eexists σ32; split => //. *)
(*       apply: has_trace_add_empty. *)
(*       apply: TraceStep => //. *)
(*       by apply: TraceEnd. *)
(*   - move => [σ11 σ21] σ31 σ32 e Hinv /(Hmstep3 _ _ _ Hinv) [σ12 [σ22 [? ?]]]. *)
(*     eexists (σ12, σ22). split => //. *)
(*     apply: has_trace_add_empty. *)
(*     apply: TraceStep => //. *)
(*     by apply: TraceEnd. *)
(* Qed. *)

Definition next_states {EV} (m : module EV) (σ : m.(m_state)) : propset (option (event EV) * m.(m_state)) :=
  {[ eσ | ∃ e, Vis <$> e = eσ.1 ∧ m.(m_step) σ e eσ.2 ]} ∪ {[ eσ | m.(m_is_ub) σ ]}.

Lemma in_next_states_has_trace {EV} (m : module EV) e σ1 σ2 :
  (e, σ2) ∈ next_states m σ1 → σ1 ~{ m, option_list e }~> σ2.
Proof.
  move => [[? /= [<- ?]]| ?].
  - apply: has_trace_add_empty. apply: TraceStep => //. by apply: TraceEnd.
  - by apply: TraceUb.
Qed.

Definition all_states_in {A B} (a : propset A) (e : propset B) (Φ : A → B → Prop) : Prop :=
  ∀ x, x ∈ a → ∃ y, y ∈ e ∧ Φ x y.

Definition all_states_in_equiv {A B} (a : propset A) (e : propset B) (Φ : A → B → Prop) : Prop :=
  all_states_in a e Φ ∧ all_states_in e a (flip Φ).

Global Instance all_states_in_proper {A B} : Proper ((≡) ==> (≡) ==> (pointwise_relation A (pointwise_relation B impl)) ==> impl) (@all_states_in A B).
Proof.
  move => a1 a2 Ha e1 e2 He Φ1 Φ2 HΦ Hall x. rewrite -Ha => Hx.
  case: (Hall _ Hx) => y. rewrite He => -[??]. eexists. split => //.
  by apply: HΦ.
Qed.

Global Instance all_states_in_equiv_proper {A B} : Proper ((≡) ==> (≡) ==> (pointwise_relation A (pointwise_relation B impl)) ==> impl) (@all_states_in_equiv A B).
Proof.
  move => ???????? HΦ [??]. split; [ by apply: all_states_in_proper|].
  apply: all_states_in_proper; [..| done] => //. move => ?? /=?. by apply: HΦ.
Qed.

Definition deterministic_step {EV} (m : module EV) (σ1 : m.(m_state)) (e : option EV) (σ2 : m.(m_state)) : Prop :=
  m.(m_step) σ1 e σ2 ∧ (∀ e' σ2', m.(m_step) σ1 e' σ2' → e' = e ∧ σ2' = σ2).

Lemma next_states_det {EV} (m : module EV) σ1 e σ2:
  deterministic_step m σ1 e σ2 → ¬ m.(m_is_ub) σ1 →
  next_states m σ1 ≡ {[(Vis <$> e, σ2)]}.
Proof.
  move => [Hdet1 Hdet2] Hub [??]. split.
  - move => [[?/=[<- /Hdet2 ?]]|//]. naive_solver.
  - move => [<- <-]. left. set_solver.
Qed.

Lemma next_states_empty {EV} (m : module EV) σ1:
  (¬ ∃ e σ2, m.(m_step) σ1 e σ2) → ¬ m.(m_is_ub) σ1 →
  next_states m σ1 ≡ ∅.
Proof. move => Hnotstep Hub [??]. split; set_solver. Qed.

Lemma all_states_in_equiv_singleton {A B} a e x y (Φ : A → B → Prop) :
  a ≡ {[ x ]} →
  e ≡ {[ y ]} →
  Φ x y →
  all_states_in_equiv a e Φ.
Proof. move => -> -> ?. split => ?; set_solver. Qed.

Lemma all_states_in_equiv_empty {A B} a e (Φ : A → B → Prop) :
  a ≡ ∅ →
  e ≡ ∅ →
  all_states_in_equiv a e Φ.
Proof. move => -> ->. split => ?; set_solver. Qed.

Lemma next_states_implies_refines {EV} (m1 m2 : mod_state EV) (inv : m1.(m_state) → m2.(m_state) → Prop):
  inv m1.(ms_state) m2.(ms_state) →
  (∀ σi σs, inv σi σs → all_states_in (next_states m1 σi) (next_states m2 σs) (λ eσi2 eσs2,
      m2.(m_is_ub) σs ∨ (eσi2.1 = eσs2.1 ∧ (m2.(m_is_ub) eσs2.2 ∨ inv eσi2.2 eσs2.2)) )) →
  m1 ⊑ m2.
Proof.
  move => Hinvinit Hinvstep.
  constructor => // κs [σi2].
  move: m1.(ms_state) m2.(ms_state) Hinvinit => σi1 σs1 Hinv Hsteps.
  elim: Hsteps σs1 Hinv => {σi1 σi2 κs}.
  - by eauto using TraceEnd.
  - move => σi1 σi2 σi3 κ κs Hstep Hsteps IH σs1 Hinv.
    case: (Hinvstep _ _ Hinv (Vis<$> κ, σi2)). { set_solver. }
    move => [? σ2] [/in_next_states_has_trace ? /= [ Hub | [? Hor]]]; simplify_eq/=.
    { eexists _. by apply: TraceUbRefl. }
    case: Hor => [? | Hinv2]. { exists σ2. apply: has_trace_trans => //. by apply: TraceUb. }
    case: (IH _ Hinv2) => ? ?.
    eexists. by apply: has_trace_trans.
  - move => σi1 ?? ? σs Hinv.
    case: (Hinvstep _ _ Hinv (Some Ub, σi1)). { set_solver. }
    move => [? ?] [Hin [? |[??]]]; simplify_eq/=.
    { eexists _. by apply: TraceUbRefl. }
    eexists. apply: TraceUbRefl. case: Hin; [ | set_solver].
    by move => [[?|][/=??]].
Qed.

Lemma next_states_implies_refines_equiv {EV} (m1 m2 : mod_state EV) (inv : m1.(m_state) → m2.(m_state) → Prop):
  inv m1.(ms_state) m2.(ms_state) →
  (∀ σi σs, inv σi σs → all_states_in_equiv (next_states m1 σi) (next_states m2 σs) (λ eσi2 eσs2,
      (m1.(m_is_ub) σi ∧ m2.(m_is_ub) σs) ∨ (eσi2.1 = eσs2.1 ∧ ((m1.(m_is_ub) eσi2.2 ∧ m2.(m_is_ub) eσs2.2) ∨ inv eσi2.2 eσs2.2)) )) →
  refines_equiv m1 m2.
Proof.
  move => Hinvinit Hinvstep.
  split.
  - apply: (next_states_implies_refines m1 m2 inv) => // σi σs Hinv.
    case: (Hinvstep _ _ Hinv) => ? _.
    apply: all_states_in_proper => // -[? ?] [??] /= ?. naive_solver.
  - apply: (next_states_implies_refines m2 m1 (flip inv)) => // σi σs Hinv.
    case: (Hinvstep _ _ Hinv) => _ ?.
    apply: all_states_in_proper => // -[? ?] [??] /= ?. naive_solver.
Qed.

Inductive wp {EV} (m1 m2 : module EV) : nat → m1.(m_state) -> m2.(m_state) -> Prop :=
| Wp_step σi1 σs1 n:
    (* This is incomplete if the inital state is UB but that is pretty weird anyway.  *)
    ¬ m1.(m_is_ub) σi1 ∧
    (∀ σi2 κ n', n = S n' → m1.(m_step) σi1 κ σi2 -> ∃ σs2,
      σs1 ~{ m2, option_list (Vis <$> κ) ++ [Ub] }~> σs2 ∨
      (σs1 ~{ m2, option_list (Vis <$> κ) }~> σs2 ∧ wp m1 m2 n' σi2 σs2)) ->
    wp m1 m2 n σi1 σs1
.

Lemma wp_implies_refines {EV} (m1 m2 : mod_state EV):
  (∀ n, wp m1 m2 n m1.(ms_state) m2.(ms_state)) →
  m1 ⊑ m2.
Proof.
  move => Hwp.
  constructor => κs [σi].
  move: m1.(ms_state) Hwp => σi1.
  move: m2.(ms_state) => σs1.
  move => Hwp Hsteps.
  move: σs1 Hwp. apply: forall_to_ex.
  elim: Hsteps => {σi1 σi κs}.
  - move => σi1. exists 0 => σs1 Hwp. eexists. by apply: TraceEnd.
  - move => σi1 σi2 σi3 κ κs Hstep Hsteps [n IH]. exists (S n) => σs1 Hwp.
    inversion_clear Hwp as [??? [? Hwp2]]; subst.
    have [|σs2 [/has_trace_app_inv [? [? /has_trace_ub_inv [σub [? ?]]]]|[? {}Hwp]]]:= (Hwp2 _ _ n _ Hstep) => //. {
      exists σub. apply: (has_trace_trans) => //. apply: (has_trace_trans []) => //. by apply: TraceUb.
    }
    have [σend ?]:= IH _ Hwp. eexists σend.
    by apply: has_trace_trans.
  - move => σ1 ???. exists 0 => ? Hwp.
    inversion_clear Hwp. naive_solver.
Qed.

Ltac invert_all_tac f :=
  let do_invert H := inversion H; clear H in
  repeat lazymatch goal with
         | H : f |- _ => do_invert H
         | H : f _ |- _ => do_invert H
         | H : f _ _|- _ => do_invert H
         | H : f _ _ _|- _ => do_invert H
         | H : f _ _ _ _|- _ => do_invert H
         | H : f _ _ _ _ _|- _ => do_invert H
         | H : f _ _ _ _ _ _|- _ => do_invert H
         | H : f _ _ _ _ _ _ _|- _ => do_invert H
         | H : f _ _ _ _ _ _ _ _|- _ => do_invert H
         | H : f _ _ _ _ _ _ _ _ _|- _ => do_invert H
         end; simplify_eq/=.

Tactic Notation "invert_all" constr(f) := invert_all_tac f.


Ltac inv_step := invert_all @m_step.

Definition module_empty {A} : module A := {|
  m_state := unit;
  m_step _ _ _ := False;
  m_is_ub s := False;
|}.
Global Instance module_empty_inst A : Empty (module A) := module_empty.

(*** Tests *)

(*
  TODO: prove the following refinement for which wp is probably not enough

            A     B
           /- 2  --- 3
  spec: 1 -
           \- 2' --- 4
            A     C

                  B
           A     /- 3
  impl: 1 --- 2 -
                 \- 4
                 C

*)
Module test.

(*   2
  1 --- 2 (done)
 *)
Inductive mod1_step : bool → option nat → bool → Prop :=
| T1False: mod1_step false (Some 2) true.


Definition mod1 : module nat := {|
  m_state := bool;
  m_step := mod1_step;
  m_is_ub s:= False;
|}.

(*         2
  1 --- 2 --- 3 (done)
 *)
Inductive mod2_state := | S1 | S2 | S3.
Inductive mod2_step : mod2_state → option nat → mod2_state → Prop :=
| T2S1: mod2_step S1 None S2
| T2S2: mod2_step S2 (Some 2) S3.
Definition mod2 : module nat := {|
  m_state := mod2_state;
  m_step := mod2_step;
  m_is_ub s:= False;
|}.

Definition t2_to_t1_inv (σ1 : mod2_state) (σ2 : bool) : Prop :=
  σ2 = match σ1 with
  | S1 | S2 => false
  | _ => true
  end.
Lemma test_refines1 :
  MS mod2 S1 ⊑ MS mod1 false.
Proof.
  apply (inv_implies_refines (MS mod2 S1) (MS mod1 false) t2_to_t1_inv).
  - done.
  - naive_solver.
  - move => σi1 σs1 σi2 e -> ?. inv_step; eexists _; right; split => //.
    + by apply: TraceEnd.
    + apply: TraceStepSome; last by apply: TraceEnd. constructor.
Qed.

Definition mod_loop {A} : module A := {|
  m_state := unit;
  m_step _ e _ := e = None;
  m_is_ub s:= False;
|}.
Lemma test_refines2 {A} (m : mod_state A) :
  MS mod_loop tt ⊑ m.
Proof.
  apply: (inv_implies_refines (MS mod_loop tt) m (λ _ _, True)).
  - done.
  - naive_solver.
  - move => ??????. inv_step. eexists. right. split => //. apply: TraceEnd.
Qed.

Lemma test_refines2_wp {A} (m : mod_state A) :
  MS mod_loop tt ⊑ m.
Proof.
  apply: wp_implies_refines => /=.
  move => n. elim/lt_wf_ind: n => n Hloop.
  constructor. split; first naive_solver. move => [] κ n' ??.
  inv_step. eexists. right. split; [by apply: TraceEnd|]. apply Hloop.
  lia.
Qed.


(*   1
      /- 2 (done)
  1 --
      \- 3 (stuck)
     2
 *)

Inductive stuck1_state := | S1S1 | S1S2 | S1S3.
Inductive stuck1_step : stuck1_state → option nat → stuck1_state → Prop :=
| S1_1To2: stuck1_step S1S1 (Some 1) S1S2
| S1_1To3: stuck1_step S1S1 (Some 2) S1S3.
Definition mod_stuck1 : module nat := {|
  m_state := stuck1_state;
  m_step := stuck1_step;
  m_is_ub s:= s = S1S3;
|}.

Lemma test_refines_stuck1 :
  MS mod_stuck1 S1S1 ⊑ MS mod_stuck1 S1S1.
Proof.
  apply: (inv_implies_refines (MS mod_stuck1 S1S1) (MS mod_stuck1 S1S1) (λ σ1 σ2, σ1 = σ2 ∧ σ1 ≠ S1S3)).
  - done.
  - move => [] ?[??] => //.
  - move => σi1 σs1 σi2 e [-> ?] ?. inv_step.
    + (* 1 -> 2 *) eexists _. right. split => //. apply: TraceStepSome; last by apply: TraceEnd. constructor.
    + (* 1 -> 3 *)
      eexists S1S1. left. apply: TraceStepSome; [constructor|]. by constructor.
Qed.

(*   1
      /- 2 (done)
  1 --
      \- 3 ---- 4 (stuck)
     2      3
 *)

Inductive stuck2_state := | S2S1 | S2S2 | S2S3 | S2S4.
Inductive stuck2_step : stuck2_state → option nat → stuck2_state → Prop :=
| S2_1To2: stuck2_step S2S1 (Some 1) S2S2
| S2_1To3: stuck2_step S2S1 (Some 2) S2S3
| S2_3To4: stuck2_step S2S3 (Some 3) S2S4.
Definition mod_stuck2 : module nat := {|
  m_state := stuck2_state;
  m_step := stuck2_step;
  m_is_ub s:= s = S2S4;
|}.

Definition stuck2_inv (σ1 : stuck2_state) (σ2 : stuck1_state) :=
  (* We could prove an even stronger invariant with also σ1 ≠ S2S3
  since we don't need to reestablish it for a stuck source state. *)
  σ1 ≠ S2S4 ∧
  σ2 = match σ1 with | S2S1 => S1S1 | S2S2 => S1S2 | S2S3 => S1S3 | S2S4 => S1S1 end.

Lemma test_refines_stuck2 :
  MS mod_stuck2 S2S1 ⊑ MS mod_stuck1 S1S1.
Proof.
  apply: (inv_implies_refines (MS mod_stuck2 S2S1) (MS mod_stuck1 S1S1) stuck2_inv).
  - done.
  - move => [] ?[??] => //.
  - move => σi1 σs1 σi2 e [? ->] ?. inv_step.
    + (* 1 -> 2 *) eexists _. right. split => //. apply: TraceStepSome; last by constructor. constructor.
    + (* 1 -> 3 *) eexists _. right. split => //. apply: TraceStepSome; last by constructor. constructor.
    + (* 3 -> 4 *) eexists S1S2. left. by apply: TraceUb.
Qed.

Lemma test_refines_stuck2_wp :
  MS mod_stuck2 S2S1 ⊑ MS mod_stuck1 S1S1.
Proof.
  apply: wp_implies_refines => n.
  (* S2S1 *)
  constructor.
  split => // σ2 ????. inv_step.
  - (* S2S2 *)
    eexists _. right. split. {
      apply: TraceStepSome; last by constructor. constructor.
    }
    constructor.
    split => // {}σ2 ????; inv_step.
  - (* S2S3 *)
    eexists _. right. split. {
      apply: TraceStepSome; last by constructor. constructor.
    }
    constructor.
    split => // {}σ2 ????.
    eexists S1S1. left. by apply: TraceUb.
Qed.

(*   1       3
      /- 2 ---- 4 (done)
  1 --
      \- 3 (stuck)
     2
 *)

Inductive stuck3_state := | S3S1 | S3S2 | S3S3 | S3S4.
Inductive stuck3_step : stuck3_state → option nat → stuck3_state → Prop :=
| S3_1To2: stuck3_step S3S1 (Some 1) S3S2
| S3_1To3: stuck3_step S3S1 (Some 2) S3S3
| S3_2To4: stuck3_step S3S2 (Some 3) S3S4.
Definition mod_stuck3 : module nat := {|
  m_state := stuck3_state;
  m_step := stuck3_step;
  m_is_ub s:= s = S3S3;
|}.

Definition stuck3_inv (σ1 : stuck3_state) (σ2 : stuck1_state) :=
  σ1 ≠ S3S3 ∧
  σ2 = match σ1 with | S3S1 => S1S1 | S3S2 => S1S2 | S3S3 => S1S3 | S3S4 => S1S2 end.

(* The following is not provable: *)
Lemma test_refines_stuck3 :
  MS mod_stuck3 S3S1 ⊑ MS mod_stuck1 S1S1.
Proof.
  apply: (inv_implies_refines (MS mod_stuck3 S3S1) (MS mod_stuck1 S1S1) stuck3_inv).
  - done.
  - move => [] ?[??] => //.
  - move => σi1 σs1 σi2 e [? ->] ?. inv_step.
    + (* 1 -> 2 *) eexists _. right. split => //. apply: TraceStepSome; last by constructor. constructor.
    + (* 1 -> 3 *)
      eexists S1S1. left. apply: TraceStepSome; [ constructor|]. by apply: TraceUb.
    + (* 2 -> 4 *) eexists _. right. split => //. apply: TraceStepSome; last by constructor.
      (* Not provable! *)
Abort.


Record call_event : Type := {
  call_nat : nat;
}.
(*
     Call 1
  1 -------- 2
 *)

Inductive call1_step : bool → option call_event → bool → Prop :=
| C1_1To2: call1_step false (Some ({| call_nat := 1 |})) true.
Definition mod_call1 : module call_event := {|
  m_state := bool;
  m_step := call1_step;
  m_is_ub s := False;
|}.

(*
            -> Call n     1 + n
  1 (done) ---------- 2 -------- 3
 *)

Inductive call2_state := | C2S1 | C2S2 (n : nat) | C2S3.
Inductive call2_step : call2_state → option (call_event + nat) → call2_state → Prop :=
| C2_1To2 cn: call2_step C2S1 (Some (inl cn)) (C2S2 cn.(call_nat))
| C2_2To3 n: call2_step (C2S2 n) (Some (inr (1 + n))) C2S3.
Definition mod_call2 : module _ := {|
  m_state := call2_state;
  m_step := call2_step;
  m_is_ub s := False;
|}.

Inductive call_merge_rel : option call_event → option (call_event + nat) → option nat → Prop :=
| CallMergeCall ev:
    call_merge_rel (Some ev) (Some (inl ev)) None
| CallMergeOut n:
    call_merge_rel None (Some (inr n)) (Some n).

Definition call_merge_inv (σ1 : bool * call2_state * unit) (σ2 : bool) :=
  match σ1.1.1, σ1.1.2 with
  | false, C2S3 => False
  | false, C2S2 _ => False
  | _, C2S2 n => n = 1
  | _, _ => True
  end ∧ σ2 = if σ1.1.2 is C2S3 then true else false.
Lemma test_refines_call_merge :
  MS (link mod_call1 mod_call2 (stateless_mediator call_merge_rel)) (false, C2S1, tt) ⊑ MS mod1 false.
Proof.
  apply: (inv_implies_refines (MS (link mod_call1 mod_call2 (stateless_mediator call_merge_rel)) (false, C2S1, tt)) (MS mod1 _) call_merge_inv).
  - done.
  - naive_solver.
  - move => σi1 σs1 σi2 e [??] ?.
    inv_step; match goal with | H : call_merge_rel _ _ _ |- _ => inversion H; clear H end; simplify_eq/=.
    + (* mod_call2 *)
      destruct σ1 => //. simplify_eq/=.
      exists true. right. split => //.
      apply: TraceStepSome; last by constructor. constructor.
    + (* mod_call1 *)
      exists false. right. split => //. by constructor.
Qed.

Definition call_split_inv (σ1 : bool) (σ2 : bool * call2_state * unit) :=
  if σ1 then True else σ2 = (false, C2S1, tt).
Lemma test_refines_call_split :
  MS mod1 false ⊑ MS (link mod_call1 mod_call2 (stateless_mediator call_merge_rel)) (false, C2S1, tt).
Proof.
  apply: (inv_implies_refines (MS mod1 _) (MS (link mod_call1 mod_call2 (stateless_mediator call_merge_rel)) _) call_split_inv).
  - done.
  - naive_solver.
  - move => σi1 [σs1 σs2] σi2 e Hinv ?. inv_step.
    exists (true, C2S3, tt). right. split => //=.
    apply: (TraceStepNone _ (link mod_call1 mod_call2 (stateless_mediator _)) (true, C2S2 1, tt)). {
      apply: LinkStepBoth. 3: constructor. all: constructor.
    }
    apply: TraceStepSome. 2: by constructor.
    apply: LinkStepR. constructor => //. simpl. constructor.
Qed.

Lemma test_refines_call_merge_wp :
  MS (link mod_call1 mod_call2 (stateless_mediator call_merge_rel)) (false, C2S1, tt) ⊑ MS mod1 false.
Proof.
  apply: (wp_implies_refines) => n.
  constructor. split; [naive_solver|] => σi1 n' ? ? Hstep. subst.
  inv_step; match goal with | H : call_merge_rel _ _ _ |- _ => inversion H; clear H end; simplify_eq/=.
  exists false.
  right. split. by constructor.

  constructor. split; [naive_solver|] => σi1 n' ? ? Hstep. subst.
  inv_step; match goal with | H : call_merge_rel _ _ _ |- _ => inversion H; clear H end; simplify_eq/=.
  exists true.
  right. split. { apply: TraceStepSome; last by constructor. constructor. }

  constructor. split; [naive_solver|] => σi1 n' ? ? Hstep. subst.
  inv_step; match goal with | H : call_merge_rel _ _ _ |- _ => inversion H; clear H end; simplify_eq/=.
Qed.

Lemma test_refines_call_split_wp :
  MS mod1 false ⊑ MS (link mod_call1 mod_call2 (stateless_mediator call_merge_rel)) (false, C2S1, tt).
Proof.
  apply: (wp_implies_refines) => n.
  constructor. split; [naive_solver|] => σi1 n' ? ? Hstep. subst.
  inv_step.
  exists (true, C2S3, tt). right.
  split. {
    apply: (TraceStepNone _ (link mod_call1 mod_call2 (stateless_mediator _)) (true, C2S2 1, tt)). {
      apply: LinkStepBoth. 3: constructor. all: constructor.
    }
    apply: TraceStepSome. 2: by constructor.
    apply: LinkStepR. constructor => //. simpl. constructor.
  }

  constructor. split; [naive_solver|] => σi1 n' ? ? Hstep. subst.
  inv_step.
Qed.

Definition call_equiv_inv (σ1 : bool * call2_state * unit) (σ2 : bool) :=
  match σ1, σ2 with
  | (false, C2S1, _), false => True
  | (true, C2S2 n, _), false => n = 1
  | (true, C2S3, _), true => True
  | _, _ => False
  end.

Lemma test_refines_call_equiv :
  refines_equiv (MS (link mod_call1 mod_call2 (stateless_mediator call_merge_rel)) (false, C2S1, tt)) (MS mod1 false).
Proof.
  apply: (inv_implies_refines_equiv (MS (link mod_call1 mod_call2 (stateless_mediator _)) _) (MS mod1 _) call_equiv_inv).
  - done.
  - naive_solver.
  - naive_solver.
  - move => σi1 σs1 σi2 e ? ?.
    inv_step; match goal with | H : call_merge_rel _ _ _ |- _ => inversion H; clear H end; simplify_eq/=.
    + right. exists true. destruct σ1, σs1 => //. simplify_eq. split; [by left|].
      apply: TraceStepSome; last by constructor. econstructor.
    + destruct σs1 => //. right. eexists false. split; [by left|]. apply: TraceEnd.
  - move => [[σi11 σi12] ?] σs1 σi2 e ? ?. inv_step.
    destruct σi11, σi12 => //; simplify_eq.
    (* TODO: it is quite bad that we have two subproofs here while with the other methods we only have 1 *)
    + right. eexists (true, C2S3, tt). split; [by left|].
      apply: TraceStepSome. 2: by constructor.
      apply: LinkStepR. constructor => //. simpl. constructor.
    + right. eexists (true, C2S3, tt). split; [by left|].
      apply: (TraceStepNone _ (link mod_call1 mod_call2 (stateless_mediator _)) (true, C2S2 1, tt)). {
        apply: LinkStepBoth. 3: constructor. all: constructor.
      }
      apply: TraceStepSome. 2: by constructor.
      apply: LinkStepR. constructor => //. simpl. constructor.
Qed.

(* Definition call_equiv_inv2 (σ1 : bool) (σ2 : call2_state) (σ3 : mod2_state) := *)
(*   match σ1, σ2, σ3 with *)
(*   | false, C2S1, S1 => True *)
(*   | true, C2S2 n, S2 => n = 1 *)
(*   | true, C2S3, S3 => True *)
(*   | _, _, _ => False *)
(*   end. *)

(* Lemma test_refines_call_equiv' : *)
(*   refines_equiv (link mod_call1 mod_call2 call_merge_rel) mod2. *)
(* Proof. *)
(*   apply: (link_merge_calls mod_call1 mod_call2 mod2 call_equiv_inv2). *)
(*   - done. *)
(*   - naive_solver. *)
(*   - move => σ1 σ2 ? Hinv ???. inv_step; destruct σ1, σ2 => //. *)
(*     + eexists true, (C2S2 1). split => //. apply: LinkStepBoth. 3: constructor. all: constructor. *)
(*     + eexists true, C2S3. simplify_eq/=. split => //. apply: LinkStepR. by constructor. simpl. constructor. *)
(*   - move => ?????????. *)
(*     inv_step; match goal with | H : call_merge_rel _ _ _ |- _ => inversion H; clear H end; simplify_eq/=. *)
(*   - move => σ1 σ2 σ3 ??????. *)
(*     inv_step; match goal with | H : call_merge_rel _ _ _ |- _ => inversion H; clear H end; simplify_eq/=. *)
(*     destruct σ1, σ3 => //. simplify_eq/=. exists S3. split => //. constructor. *)
(*   - move => σ1 σ2 σ3 ?????????. *)
(*     match goal with | H : call_merge_rel _ _ _ |- _ => inversion H; clear H end; simplify_eq/=. *)
(*     match goal with | H : call1_step _ _ _ |- _ => inversion H; clear H end; simplify_eq/=. *)
(*     match goal with | H : call2_step _ _ _ |- _ => inversion H; clear H end; simplify_eq/=. *)
(*     destruct σ3 => //. eexists S2. split => //. constructor. *)
(* Qed. *)

Definition call_equiv_inv2 (σ1 : bool * call2_state * unit) (σ2 : mod2_state) :=
  match σ1, σ2 with
  | (false, C2S1, _), S1 => True
  | (true, C2S2 n, _), S2 => n = 1
  | (true, C2S3, _), S3 => True
  | _, _ => False
  end.

Local Ltac solve_refines_call_next_equiv_det :=
  split; [ by repeat econstructor | move => ???; invert_all @m_step; destruct_hyps; by invert_all call_merge_rel].
Lemma test_refines_call_next_equiv :
  refines_equiv (MS (link mod_call1 mod_call2 (stateless_mediator call_merge_rel)) (false, C2S1, tt)) (MS mod2 S1).
Proof.
  apply (next_states_implies_refines_equiv (MS (link mod_call1 mod_call2 (stateless_mediator call_merge_rel)) _) (MS mod2 _) (call_equiv_inv2)).
  - done.
  - move => [[σi1 σi2] []] σs /=.
    destruct σi1, σi2, σs => //= [->|_|_].
    + apply: all_states_in_equiv_singleton;
        [ rewrite next_states_det; [done| solve_refines_call_next_equiv_det |naive_solver].. |].
      naive_solver.
    + apply: all_states_in_equiv_empty;
        (rewrite next_states_empty; [done | move => [?[??]]; inv_step | naive_solver]).
    + apply: all_states_in_equiv_singleton;
        [ rewrite next_states_det; [done| solve_refines_call_next_equiv_det |naive_solver].. |].
      naive_solver.
Qed.


End test.
